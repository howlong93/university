module sec_approx (
    //INPUT
    signed,
    //OUTPUT
)