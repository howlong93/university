module reciprocal_sqrt_rom(KEY, VALUE);
  input [14:0] KEY;
  output reg [18:0] VALUE;

  always @(KEY)begin
    case (KEY)
      15'b000_000000000001 : VALUE=19'b0111111_111111111111;
      15'b000_000000000010 : VALUE=19'b0101101_010000010100;
      15'b000_000000000011 : VALUE=19'b0100100_111100110101;
      15'b000_000000000100 : VALUE=19'b0100000_000000000000;
      15'b000_000000000101 : VALUE=19'b0011100_100111110010;
      15'b000_000000000110 : VALUE=19'b0011010_001000001100;
      15'b000_000000000111 : VALUE=19'b0011000_001100001001;
      15'b000_000000001000 : VALUE=19'b0010110_101000001010;
      15'b000_000000001001 : VALUE=19'b0010101_010101010101;
      15'b000_000000001010 : VALUE=19'b0010100_001111010001;
      15'b000_000000001011 : VALUE=19'b0010011_010010111111;
      15'b000_000000001100 : VALUE=19'b0010010_011110011010;
      15'b000_000000001101 : VALUE=19'b0010001_110000000010;
      15'b000_000000001110 : VALUE=19'b0010001_000110101101;
      15'b000_000000001111 : VALUE=19'b0010000_100001100101;
      15'b000_000000010000 : VALUE=19'b0010000_000000000000;
      15'b000_000000010001 : VALUE=19'b0001111_100001011011;
      15'b000_000000010010 : VALUE=19'b0001111_000101011100;
      15'b000_000000010011 : VALUE=19'b0001110_101011101100;
      15'b000_000000010100 : VALUE=19'b0001110_010011111001;
      15'b000_000000010101 : VALUE=19'b0001101_111101110101;
      15'b000_000000010110 : VALUE=19'b0001101_101001010001;
      15'b000_000000010111 : VALUE=19'b0001101_010110000101;
      15'b000_000000011000 : VALUE=19'b0001101_000100000110;
      15'b000_000000011001 : VALUE=19'b0001100_110011001101;
      15'b000_000000011010 : VALUE=19'b0001100_100011010011;
      15'b000_000000011011 : VALUE=19'b0001100_010100010010;
      15'b000_000000011100 : VALUE=19'b0001100_000110000101;
      15'b000_000000011101 : VALUE=19'b0001011_111000100111;
      15'b000_000000011110 : VALUE=19'b0001011_101011110101;
      15'b000_000000011111 : VALUE=19'b0001011_011111101010;
      15'b000_000000100000 : VALUE=19'b0001011_010100000101;
      15'b000_000000100001 : VALUE=19'b0001011_001001000001;
      15'b000_000000100010 : VALUE=19'b0001010_111110011101;
      15'b000_000000100011 : VALUE=19'b0001010_110100010110;
      15'b000_000000100100 : VALUE=19'b0001010_101010101011;
      15'b000_000000100101 : VALUE=19'b0001010_100001011000;
      15'b000_000000100110 : VALUE=19'b0001010_011000011101;
      15'b000_000000100111 : VALUE=19'b0001010_001111111001;
      15'b000_000000101000 : VALUE=19'b0001010_000111101001;
      15'b000_000000101001 : VALUE=19'b0001001_111111101100;
      15'b000_000000101010 : VALUE=19'b0001001_111000000010;
      15'b000_000000101011 : VALUE=19'b0001001_110000101001;
      15'b000_000000101100 : VALUE=19'b0001001_101001100000;
      15'b000_000000101101 : VALUE=19'b0001001_100010100110;
      15'b000_000000101110 : VALUE=19'b0001001_011011111011;
      15'b000_000000101111 : VALUE=19'b0001001_010101011110;
      15'b000_000000110000 : VALUE=19'b0001001_001111001101;
      15'b000_000000110001 : VALUE=19'b0001001_001001001001;
      15'b000_000000110010 : VALUE=19'b0001001_000011010001;
      15'b000_000000110011 : VALUE=19'b0001000_111101100100;
      15'b000_000000110100 : VALUE=19'b0001000_111000000001;
      15'b000_000000110101 : VALUE=19'b0001000_110010101000;
      15'b000_000000110110 : VALUE=19'b0001000_101101011001;
      15'b000_000000110111 : VALUE=19'b0001000_101000010011;
      15'b000_000000111000 : VALUE=19'b0001000_100011010110;
      15'b000_000000111001 : VALUE=19'b0001000_011110100010;
      15'b000_000000111010 : VALUE=19'b0001000_011001110101;
      15'b000_000000111011 : VALUE=19'b0001000_010101010000;
      15'b000_000000111100 : VALUE=19'b0001000_010000110011;
      15'b000_000000111101 : VALUE=19'b0001000_001100011100;
      15'b000_000000111110 : VALUE=19'b0001000_001000001100;
      15'b000_000000111111 : VALUE=19'b0001000_000100000011;
      15'b000_000001000000 : VALUE=19'b0001000_000000000000;
      15'b000_000001000001 : VALUE=19'b0000111_111100000011;
      15'b000_000001000010 : VALUE=19'b0000111_111000001100;
      15'b000_000001000011 : VALUE=19'b0000111_110100011010;
      15'b000_000001000100 : VALUE=19'b0000111_110000101110;
      15'b000_000001000101 : VALUE=19'b0000111_101101000110;
      15'b000_000001000110 : VALUE=19'b0000111_101001100100;
      15'b000_000001000111 : VALUE=19'b0000111_100110000111;
      15'b000_000001001000 : VALUE=19'b0000111_100010101110;
      15'b000_000001001001 : VALUE=19'b0000111_011111011010;
      15'b000_000001001010 : VALUE=19'b0000111_011100001010;
      15'b000_000001001011 : VALUE=19'b0000111_011000111110;
      15'b000_000001001100 : VALUE=19'b0000111_010101110110;
      15'b000_000001001101 : VALUE=19'b0000111_010010110010;
      15'b000_000001001110 : VALUE=19'b0000111_001111110010;
      15'b000_000001001111 : VALUE=19'b0000111_001100110110;
      15'b000_000001010000 : VALUE=19'b0000111_001001111101;
      15'b000_000001010001 : VALUE=19'b0000111_000111000111;
      15'b000_000001010010 : VALUE=19'b0000111_000100010101;
      15'b000_000001010011 : VALUE=19'b0000111_000001100110;
      15'b000_000001010100 : VALUE=19'b0000110_111110111010;
      15'b000_000001010101 : VALUE=19'b0000110_111100010010;
      15'b000_000001010110 : VALUE=19'b0000110_111001101100;
      15'b000_000001010111 : VALUE=19'b0000110_110111001001;
      15'b000_000001011000 : VALUE=19'b0000110_110100101001;
      15'b000_000001011001 : VALUE=19'b0000110_110010001011;
      15'b000_000001011010 : VALUE=19'b0000110_101111110000;
      15'b000_000001011011 : VALUE=19'b0000110_101101011000;
      15'b000_000001011100 : VALUE=19'b0000110_101011000010;
      15'b000_000001011101 : VALUE=19'b0000110_101000101111;
      15'b000_000001011110 : VALUE=19'b0000110_100110011110;
      15'b000_000001011111 : VALUE=19'b0000110_100100001111;
      15'b000_000001100000 : VALUE=19'b0000110_100010000011;
      15'b000_000001100001 : VALUE=19'b0000110_011111111001;
      15'b000_000001100010 : VALUE=19'b0000110_011101110001;
      15'b000_000001100011 : VALUE=19'b0000110_011011101010;
      15'b000_000001100100 : VALUE=19'b0000110_011001100110;
      15'b000_000001100101 : VALUE=19'b0000110_010111100100;
      15'b000_000001100110 : VALUE=19'b0000110_010101100100;
      15'b000_000001100111 : VALUE=19'b0000110_010011100110;
      15'b000_000001101000 : VALUE=19'b0000110_010001101001;
      15'b000_000001101001 : VALUE=19'b0000110_001111101111;
      15'b000_000001101010 : VALUE=19'b0000110_001101110110;
      15'b000_000001101011 : VALUE=19'b0000110_001011111110;
      15'b000_000001101100 : VALUE=19'b0000110_001010001001;
      15'b000_000001101101 : VALUE=19'b0000110_001000010101;
      15'b000_000001101110 : VALUE=19'b0000110_000110100010;
      15'b000_000001101111 : VALUE=19'b0000110_000100110010;
      15'b000_000001110000 : VALUE=19'b0000110_000011000010;
      15'b000_000001110001 : VALUE=19'b0000110_000001010100;
      15'b000_000001110010 : VALUE=19'b0000101_111111101000;
      15'b000_000001110011 : VALUE=19'b0000101_111101111101;
      15'b000_000001110100 : VALUE=19'b0000101_111100010011;
      15'b000_000001110101 : VALUE=19'b0000101_111010101011;
      15'b000_000001110110 : VALUE=19'b0000101_111001000100;
      15'b000_000001110111 : VALUE=19'b0000101_110111011111;
      15'b000_000001111000 : VALUE=19'b0000101_110101111010;
      15'b000_000001111001 : VALUE=19'b0000101_110100010111;
      15'b000_000001111010 : VALUE=19'b0000101_110010110101;
      15'b000_000001111011 : VALUE=19'b0000101_110001010101;
      15'b000_000001111100 : VALUE=19'b0000101_101111110101;
      15'b000_000001111101 : VALUE=19'b0000101_101110010111;
      15'b000_000001111110 : VALUE=19'b0000101_101100111010;
      15'b000_000001111111 : VALUE=19'b0000101_101011011110;
      15'b000_000010000000 : VALUE=19'b0000101_101010000010;
      15'b000_000010000001 : VALUE=19'b0000101_101000101000;
      15'b000_000010000010 : VALUE=19'b0000101_100111010000;
      15'b000_000010000011 : VALUE=19'b0000101_100101111000;
      15'b000_000010000100 : VALUE=19'b0000101_100100100001;
      15'b000_000010000101 : VALUE=19'b0000101_100011001011;
      15'b000_000010000110 : VALUE=19'b0000101_100001110110;
      15'b000_000010000111 : VALUE=19'b0000101_100000100010;
      15'b000_000010001000 : VALUE=19'b0000101_011111001111;
      15'b000_000010001001 : VALUE=19'b0000101_011101111100;
      15'b000_000010001010 : VALUE=19'b0000101_011100101011;
      15'b000_000010001011 : VALUE=19'b0000101_011011011011;
      15'b000_000010001100 : VALUE=19'b0000101_011010001011;
      15'b000_000010001101 : VALUE=19'b0000101_011000111101;
      15'b000_000010001110 : VALUE=19'b0000101_010111101111;
      15'b000_000010001111 : VALUE=19'b0000101_010110100010;
      15'b000_000010010000 : VALUE=19'b0000101_010101010101;
      15'b000_000010010001 : VALUE=19'b0000101_010100001010;
      15'b000_000010010010 : VALUE=19'b0000101_010010111111;
      15'b000_000010010011 : VALUE=19'b0000101_010001110101;
      15'b000_000010010100 : VALUE=19'b0000101_010000101100;
      15'b000_000010010101 : VALUE=19'b0000101_001111100100;
      15'b000_000010010110 : VALUE=19'b0000101_001110011100;
      15'b000_000010010111 : VALUE=19'b0000101_001101010101;
      15'b000_000010011000 : VALUE=19'b0000101_001100001111;
      15'b000_000010011001 : VALUE=19'b0000101_001011001001;
      15'b000_000010011010 : VALUE=19'b0000101_001010000100;
      15'b000_000010011011 : VALUE=19'b0000101_001001000000;
      15'b000_000010011100 : VALUE=19'b0000101_000111111100;
      15'b000_000010011101 : VALUE=19'b0000101_000110111001;
      15'b000_000010011110 : VALUE=19'b0000101_000101110111;
      15'b000_000010011111 : VALUE=19'b0000101_000100110101;
      15'b000_000010100000 : VALUE=19'b0000101_000011110100;
      15'b000_000010100001 : VALUE=19'b0000101_000010110100;
      15'b000_000010100010 : VALUE=19'b0000101_000001110100;
      15'b000_000010100011 : VALUE=19'b0000101_000000110101;
      15'b000_000010100100 : VALUE=19'b0000100_111111110110;
      15'b000_000010100101 : VALUE=19'b0000100_111110111000;
      15'b000_000010100110 : VALUE=19'b0000100_111101111010;
      15'b000_000010100111 : VALUE=19'b0000100_111100111101;
      15'b000_000010101000 : VALUE=19'b0000100_111100000001;
      15'b000_000010101001 : VALUE=19'b0000100_111011000101;
      15'b000_000010101010 : VALUE=19'b0000100_111010001010;
      15'b000_000010101011 : VALUE=19'b0000100_111001001111;
      15'b000_000010101100 : VALUE=19'b0000100_111000010100;
      15'b000_000010101101 : VALUE=19'b0000100_110111011010;
      15'b000_000010101110 : VALUE=19'b0000100_110110100001;
      15'b000_000010101111 : VALUE=19'b0000100_110101101000;
      15'b000_000010110000 : VALUE=19'b0000100_110100110000;
      15'b000_000010110001 : VALUE=19'b0000100_110011111000;
      15'b000_000010110010 : VALUE=19'b0000100_110011000001;
      15'b000_000010110011 : VALUE=19'b0000100_110010001010;
      15'b000_000010110100 : VALUE=19'b0000100_110001010011;
      15'b000_000010110101 : VALUE=19'b0000100_110000011101;
      15'b000_000010110110 : VALUE=19'b0000100_101111100111;
      15'b000_000010110111 : VALUE=19'b0000100_101110110010;
      15'b000_000010111000 : VALUE=19'b0000100_101101111110;
      15'b000_000010111001 : VALUE=19'b0000100_101101001001;
      15'b000_000010111010 : VALUE=19'b0000100_101100010101;
      15'b000_000010111011 : VALUE=19'b0000100_101011100010;
      15'b000_000010111100 : VALUE=19'b0000100_101010101111;
      15'b000_000010111101 : VALUE=19'b0000100_101001111100;
      15'b000_000010111110 : VALUE=19'b0000100_101001001010;
      15'b000_000010111111 : VALUE=19'b0000100_101000011000;
      15'b000_000011000000 : VALUE=19'b0000100_100111100111;
      15'b000_000011000001 : VALUE=19'b0000100_100110110110;
      15'b000_000011000010 : VALUE=19'b0000100_100110000101;
      15'b000_000011000011 : VALUE=19'b0000100_100101010101;
      15'b000_000011000100 : VALUE=19'b0000100_100100100101;
      15'b000_000011000101 : VALUE=19'b0000100_100011110101;
      15'b000_000011000110 : VALUE=19'b0000100_100011000110;
      15'b000_000011000111 : VALUE=19'b0000100_100010010111;
      15'b000_000011001000 : VALUE=19'b0000100_100001101000;
      15'b000_000011001001 : VALUE=19'b0000100_100000111010;
      15'b000_000011001010 : VALUE=19'b0000100_100000001100;
      15'b000_000011001011 : VALUE=19'b0000100_011111011111;
      15'b000_000011001100 : VALUE=19'b0000100_011110110010;
      15'b000_000011001101 : VALUE=19'b0000100_011110000101;
      15'b000_000011001110 : VALUE=19'b0000100_011101011000;
      15'b000_000011001111 : VALUE=19'b0000100_011100101100;
      15'b000_000011010000 : VALUE=19'b0000100_011100000000;
      15'b000_000011010001 : VALUE=19'b0000100_011011010101;
      15'b000_000011010010 : VALUE=19'b0000100_011010101010;
      15'b000_000011010011 : VALUE=19'b0000100_011001111111;
      15'b000_000011010100 : VALUE=19'b0000100_011001010100;
      15'b000_000011010101 : VALUE=19'b0000100_011000101010;
      15'b000_000011010110 : VALUE=19'b0000100_011000000000;
      15'b000_000011010111 : VALUE=19'b0000100_010111010110;
      15'b000_000011011000 : VALUE=19'b0000100_010110101101;
      15'b000_000011011001 : VALUE=19'b0000100_010110000011;
      15'b000_000011011010 : VALUE=19'b0000100_010101011011;
      15'b000_000011011011 : VALUE=19'b0000100_010100110010;
      15'b000_000011011100 : VALUE=19'b0000100_010100001010;
      15'b000_000011011101 : VALUE=19'b0000100_010011100010;
      15'b000_000011011110 : VALUE=19'b0000100_010010111010;
      15'b000_000011011111 : VALUE=19'b0000100_010010010010;
      15'b000_000011100000 : VALUE=19'b0000100_010001101011;
      15'b000_000011100001 : VALUE=19'b0000100_010001000100;
      15'b000_000011100010 : VALUE=19'b0000100_010000011110;
      15'b000_000011100011 : VALUE=19'b0000100_001111110111;
      15'b000_000011100100 : VALUE=19'b0000100_001111010001;
      15'b000_000011100101 : VALUE=19'b0000100_001110101011;
      15'b000_000011100110 : VALUE=19'b0000100_001110000101;
      15'b000_000011100111 : VALUE=19'b0000100_001101100000;
      15'b000_000011101000 : VALUE=19'b0000100_001100111011;
      15'b000_000011101001 : VALUE=19'b0000100_001100010110;
      15'b000_000011101010 : VALUE=19'b0000100_001011110001;
      15'b000_000011101011 : VALUE=19'b0000100_001011001100;
      15'b000_000011101100 : VALUE=19'b0000100_001010101000;
      15'b000_000011101101 : VALUE=19'b0000100_001010000100;
      15'b000_000011101110 : VALUE=19'b0000100_001001100000;
      15'b000_000011101111 : VALUE=19'b0000100_001000111101;
      15'b000_000011110000 : VALUE=19'b0000100_001000011001;
      15'b000_000011110001 : VALUE=19'b0000100_000111110110;
      15'b000_000011110010 : VALUE=19'b0000100_000111010011;
      15'b000_000011110011 : VALUE=19'b0000100_000110110001;
      15'b000_000011110100 : VALUE=19'b0000100_000110001110;
      15'b000_000011110101 : VALUE=19'b0000100_000101101100;
      15'b000_000011110110 : VALUE=19'b0000100_000101001010;
      15'b000_000011110111 : VALUE=19'b0000100_000100101000;
      15'b000_000011111000 : VALUE=19'b0000100_000100000110;
      15'b000_000011111001 : VALUE=19'b0000100_000011100101;
      15'b000_000011111010 : VALUE=19'b0000100_000011000011;
      15'b000_000011111011 : VALUE=19'b0000100_000010100010;
      15'b000_000011111100 : VALUE=19'b0000100_000010000010;
      15'b000_000011111101 : VALUE=19'b0000100_000001100001;
      15'b000_000011111110 : VALUE=19'b0000100_000001000000;
      15'b000_000011111111 : VALUE=19'b0000100_000000100000;
      15'b000_000100000000 : VALUE=19'b0000100_000000000000;
      15'b000_000100000001 : VALUE=19'b0000011_111111100000;
      15'b000_000100000010 : VALUE=19'b0000011_111111000000;
      15'b000_000100000011 : VALUE=19'b0000011_111110100001;
      15'b000_000100000100 : VALUE=19'b0000011_111110000001;
      15'b000_000100000101 : VALUE=19'b0000011_111101100010;
      15'b000_000100000110 : VALUE=19'b0000011_111101000011;
      15'b000_000100000111 : VALUE=19'b0000011_111100100100;
      15'b000_000100001000 : VALUE=19'b0000011_111100000110;
      15'b000_000100001001 : VALUE=19'b0000011_111011100111;
      15'b000_000100001010 : VALUE=19'b0000011_111011001001;
      15'b000_000100001011 : VALUE=19'b0000011_111010101011;
      15'b000_000100001100 : VALUE=19'b0000011_111010001101;
      15'b000_000100001101 : VALUE=19'b0000011_111001101111;
      15'b000_000100001110 : VALUE=19'b0000011_111001010010;
      15'b000_000100001111 : VALUE=19'b0000011_111000110100;
      15'b000_000100010000 : VALUE=19'b0000011_111000010111;
      15'b000_000100010001 : VALUE=19'b0000011_110111111010;
      15'b000_000100010010 : VALUE=19'b0000011_110111011101;
      15'b000_000100010011 : VALUE=19'b0000011_110111000000;
      15'b000_000100010100 : VALUE=19'b0000011_110110100011;
      15'b000_000100010101 : VALUE=19'b0000011_110110000111;
      15'b000_000100010110 : VALUE=19'b0000011_110101101010;
      15'b000_000100010111 : VALUE=19'b0000011_110101001110;
      15'b000_000100011000 : VALUE=19'b0000011_110100110010;
      15'b000_000100011001 : VALUE=19'b0000011_110100010110;
      15'b000_000100011010 : VALUE=19'b0000011_110011111010;
      15'b000_000100011011 : VALUE=19'b0000011_110011011111;
      15'b000_000100011100 : VALUE=19'b0000011_110011000011;
      15'b000_000100011101 : VALUE=19'b0000011_110010101000;
      15'b000_000100011110 : VALUE=19'b0000011_110010001101;
      15'b000_000100011111 : VALUE=19'b0000011_110001110010;
      15'b000_000100100000 : VALUE=19'b0000011_110001010111;
      15'b000_000100100001 : VALUE=19'b0000011_110000111100;
      15'b000_000100100010 : VALUE=19'b0000011_110000100010;
      15'b000_000100100011 : VALUE=19'b0000011_110000000111;
      15'b000_000100100100 : VALUE=19'b0000011_101111101101;
      15'b000_000100100101 : VALUE=19'b0000011_101111010011;
      15'b000_000100100110 : VALUE=19'b0000011_101110111001;
      15'b000_000100100111 : VALUE=19'b0000011_101110011111;
      15'b000_000100101000 : VALUE=19'b0000011_101110000101;
      15'b000_000100101001 : VALUE=19'b0000011_101101101011;
      15'b000_000100101010 : VALUE=19'b0000011_101101010010;
      15'b000_000100101011 : VALUE=19'b0000011_101100111000;
      15'b000_000100101100 : VALUE=19'b0000011_101100011111;
      15'b000_000100101101 : VALUE=19'b0000011_101100000110;
      15'b000_000100101110 : VALUE=19'b0000011_101011101101;
      15'b000_000100101111 : VALUE=19'b0000011_101011010100;
      15'b000_000100110000 : VALUE=19'b0000011_101010111011;
      15'b000_000100110001 : VALUE=19'b0000011_101010100010;
      15'b000_000100110010 : VALUE=19'b0000011_101010001010;
      15'b000_000100110011 : VALUE=19'b0000011_101001110001;
      15'b000_000100110100 : VALUE=19'b0000011_101001011001;
      15'b000_000100110101 : VALUE=19'b0000011_101001000001;
      15'b000_000100110110 : VALUE=19'b0000011_101000101001;
      15'b000_000100110111 : VALUE=19'b0000011_101000010001;
      15'b000_000100111000 : VALUE=19'b0000011_100111111001;
      15'b000_000100111001 : VALUE=19'b0000011_100111100001;
      15'b000_000100111010 : VALUE=19'b0000011_100111001010;
      15'b000_000100111011 : VALUE=19'b0000011_100110110010;
      15'b000_000100111100 : VALUE=19'b0000011_100110011011;
      15'b000_000100111101 : VALUE=19'b0000011_100110000011;
      15'b000_000100111110 : VALUE=19'b0000011_100101101100;
      15'b000_000100111111 : VALUE=19'b0000011_100101010101;
      15'b000_000101000000 : VALUE=19'b0000011_100100111110;
      15'b000_000101000001 : VALUE=19'b0000011_100100100111;
      15'b000_000101000010 : VALUE=19'b0000011_100100010001;
      15'b000_000101000011 : VALUE=19'b0000011_100011111010;
      15'b000_000101000100 : VALUE=19'b0000011_100011100100;
      15'b000_000101000101 : VALUE=19'b0000011_100011001101;
      15'b000_000101000110 : VALUE=19'b0000011_100010110111;
      15'b000_000101000111 : VALUE=19'b0000011_100010100001;
      15'b000_000101001000 : VALUE=19'b0000011_100010001010;
      15'b000_000101001001 : VALUE=19'b0000011_100001110100;
      15'b000_000101001010 : VALUE=19'b0000011_100001011111;
      15'b000_000101001011 : VALUE=19'b0000011_100001001001;
      15'b000_000101001100 : VALUE=19'b0000011_100000110011;
      15'b000_000101001101 : VALUE=19'b0000011_100000011101;
      15'b000_000101001110 : VALUE=19'b0000011_100000001000;
      15'b000_000101001111 : VALUE=19'b0000011_011111110010;
      15'b000_000101010000 : VALUE=19'b0000011_011111011101;
      15'b000_000101010001 : VALUE=19'b0000011_011111001000;
      15'b000_000101010010 : VALUE=19'b0000011_011110110011;
      15'b000_000101010011 : VALUE=19'b0000011_011110011110;
      15'b000_000101010100 : VALUE=19'b0000011_011110001001;
      15'b000_000101010101 : VALUE=19'b0000011_011101110100;
      15'b000_000101010110 : VALUE=19'b0000011_011101011111;
      15'b000_000101010111 : VALUE=19'b0000011_011101001010;
      15'b000_000101011000 : VALUE=19'b0000011_011100110110;
      15'b000_000101011001 : VALUE=19'b0000011_011100100001;
      15'b000_000101011010 : VALUE=19'b0000011_011100001101;
      15'b000_000101011011 : VALUE=19'b0000011_011011111001;
      15'b000_000101011100 : VALUE=19'b0000011_011011100100;
      15'b000_000101011101 : VALUE=19'b0000011_011011010000;
      15'b000_000101011110 : VALUE=19'b0000011_011010111100;
      15'b000_000101011111 : VALUE=19'b0000011_011010101000;
      15'b000_000101100000 : VALUE=19'b0000011_011010010100;
      15'b000_000101100001 : VALUE=19'b0000011_011010000001;
      15'b000_000101100010 : VALUE=19'b0000011_011001101101;
      15'b000_000101100011 : VALUE=19'b0000011_011001011001;
      15'b000_000101100100 : VALUE=19'b0000011_011001000110;
      15'b000_000101100101 : VALUE=19'b0000011_011000110010;
      15'b000_000101100110 : VALUE=19'b0000011_011000011111;
      15'b000_000101100111 : VALUE=19'b0000011_011000001011;
      15'b000_000101101000 : VALUE=19'b0000011_010111111000;
      15'b000_000101101001 : VALUE=19'b0000011_010111100101;
      15'b000_000101101010 : VALUE=19'b0000011_010111010010;
      15'b000_000101101011 : VALUE=19'b0000011_010110111111;
      15'b000_000101101100 : VALUE=19'b0000011_010110101100;
      15'b000_000101101101 : VALUE=19'b0000011_010110011001;
      15'b000_000101101110 : VALUE=19'b0000011_010110000110;
      15'b000_000101101111 : VALUE=19'b0000011_010101110100;
      15'b000_000101110000 : VALUE=19'b0000011_010101100001;
      15'b000_000101110001 : VALUE=19'b0000011_010101001111;
      15'b000_000101110010 : VALUE=19'b0000011_010100111100;
      15'b000_000101110011 : VALUE=19'b0000011_010100101010;
      15'b000_000101110100 : VALUE=19'b0000011_010100011000;
      15'b000_000101110101 : VALUE=19'b0000011_010100000101;
      15'b000_000101110110 : VALUE=19'b0000011_010011110011;
      15'b000_000101110111 : VALUE=19'b0000011_010011100001;
      15'b000_000101111000 : VALUE=19'b0000011_010011001111;
      15'b000_000101111001 : VALUE=19'b0000011_010010111101;
      15'b000_000101111010 : VALUE=19'b0000011_010010101011;
      15'b000_000101111011 : VALUE=19'b0000011_010010011001;
      15'b000_000101111100 : VALUE=19'b0000011_010010001000;
      15'b000_000101111101 : VALUE=19'b0000011_010001110110;
      15'b000_000101111110 : VALUE=19'b0000011_010001100100;
      15'b000_000101111111 : VALUE=19'b0000011_010001010011;
      15'b000_000110000000 : VALUE=19'b0000011_010001000001;
      15'b000_000110000001 : VALUE=19'b0000011_010000110000;
      15'b000_000110000010 : VALUE=19'b0000011_010000011111;
      15'b000_000110000011 : VALUE=19'b0000011_010000001110;
      15'b000_000110000100 : VALUE=19'b0000011_001111111100;
      15'b000_000110000101 : VALUE=19'b0000011_001111101011;
      15'b000_000110000110 : VALUE=19'b0000011_001111011010;
      15'b000_000110000111 : VALUE=19'b0000011_001111001001;
      15'b000_000110001000 : VALUE=19'b0000011_001110111000;
      15'b000_000110001001 : VALUE=19'b0000011_001110100111;
      15'b000_000110001010 : VALUE=19'b0000011_001110010111;
      15'b000_000110001011 : VALUE=19'b0000011_001110000110;
      15'b000_000110001100 : VALUE=19'b0000011_001101110101;
      15'b000_000110001101 : VALUE=19'b0000011_001101100101;
      15'b000_000110001110 : VALUE=19'b0000011_001101010100;
      15'b000_000110001111 : VALUE=19'b0000011_001101000100;
      15'b000_000110010000 : VALUE=19'b0000011_001100110011;
      15'b000_000110010001 : VALUE=19'b0000011_001100100011;
      15'b000_000110010010 : VALUE=19'b0000011_001100010011;
      15'b000_000110010011 : VALUE=19'b0000011_001100000010;
      15'b000_000110010100 : VALUE=19'b0000011_001011110010;
      15'b000_000110010101 : VALUE=19'b0000011_001011100010;
      15'b000_000110010110 : VALUE=19'b0000011_001011010010;
      15'b000_000110010111 : VALUE=19'b0000011_001011000010;
      15'b000_000110011000 : VALUE=19'b0000011_001010110010;
      15'b000_000110011001 : VALUE=19'b0000011_001010100010;
      15'b000_000110011010 : VALUE=19'b0000011_001010010010;
      15'b000_000110011011 : VALUE=19'b0000011_001010000011;
      15'b000_000110011100 : VALUE=19'b0000011_001001110011;
      15'b000_000110011101 : VALUE=19'b0000011_001001100011;
      15'b000_000110011110 : VALUE=19'b0000011_001001010100;
      15'b000_000110011111 : VALUE=19'b0000011_001001000100;
      15'b000_000110100000 : VALUE=19'b0000011_001000110101;
      15'b000_000110100001 : VALUE=19'b0000011_001000100101;
      15'b000_000110100010 : VALUE=19'b0000011_001000010110;
      15'b000_000110100011 : VALUE=19'b0000011_001000000111;
      15'b000_000110100100 : VALUE=19'b0000011_000111110111;
      15'b000_000110100101 : VALUE=19'b0000011_000111101000;
      15'b000_000110100110 : VALUE=19'b0000011_000111011001;
      15'b000_000110100111 : VALUE=19'b0000011_000111001010;
      15'b000_000110101000 : VALUE=19'b0000011_000110111011;
      15'b000_000110101001 : VALUE=19'b0000011_000110101100;
      15'b000_000110101010 : VALUE=19'b0000011_000110011101;
      15'b000_000110101011 : VALUE=19'b0000011_000110001110;
      15'b000_000110101100 : VALUE=19'b0000011_000101111111;
      15'b000_000110101101 : VALUE=19'b0000011_000101110000;
      15'b000_000110101110 : VALUE=19'b0000011_000101100010;
      15'b000_000110101111 : VALUE=19'b0000011_000101010011;
      15'b000_000110110000 : VALUE=19'b0000011_000101000100;
      15'b000_000110110001 : VALUE=19'b0000011_000100110110;
      15'b000_000110110010 : VALUE=19'b0000011_000100100111;
      15'b000_000110110011 : VALUE=19'b0000011_000100011001;
      15'b000_000110110100 : VALUE=19'b0000011_000100001010;
      15'b000_000110110101 : VALUE=19'b0000011_000011111100;
      15'b000_000110110110 : VALUE=19'b0000011_000011101110;
      15'b000_000110110111 : VALUE=19'b0000011_000011011111;
      15'b000_000110111000 : VALUE=19'b0000011_000011010001;
      15'b000_000110111001 : VALUE=19'b0000011_000011000011;
      15'b000_000110111010 : VALUE=19'b0000011_000010110101;
      15'b000_000110111011 : VALUE=19'b0000011_000010100111;
      15'b000_000110111100 : VALUE=19'b0000011_000010011001;
      15'b000_000110111101 : VALUE=19'b0000011_000010001011;
      15'b000_000110111110 : VALUE=19'b0000011_000001111101;
      15'b000_000110111111 : VALUE=19'b0000011_000001101111;
      15'b000_000111000000 : VALUE=19'b0000011_000001100001;
      15'b000_000111000001 : VALUE=19'b0000011_000001010011;
      15'b000_000111000010 : VALUE=19'b0000011_000001000110;
      15'b000_000111000011 : VALUE=19'b0000011_000000111000;
      15'b000_000111000100 : VALUE=19'b0000011_000000101010;
      15'b000_000111000101 : VALUE=19'b0000011_000000011101;
      15'b000_000111000110 : VALUE=19'b0000011_000000001111;
      15'b000_000111000111 : VALUE=19'b0000011_000000000010;
      15'b000_000111001000 : VALUE=19'b0000010_111111110100;
      15'b000_000111001001 : VALUE=19'b0000010_111111100111;
      15'b000_000111001010 : VALUE=19'b0000010_111111011001;
      15'b000_000111001011 : VALUE=19'b0000010_111111001100;
      15'b000_000111001100 : VALUE=19'b0000010_111110111111;
      15'b000_000111001101 : VALUE=19'b0000010_111110110001;
      15'b000_000111001110 : VALUE=19'b0000010_111110100100;
      15'b000_000111001111 : VALUE=19'b0000010_111110010111;
      15'b000_000111010000 : VALUE=19'b0000010_111110001010;
      15'b000_000111010001 : VALUE=19'b0000010_111101111101;
      15'b000_000111010010 : VALUE=19'b0000010_111101110000;
      15'b000_000111010011 : VALUE=19'b0000010_111101100011;
      15'b000_000111010100 : VALUE=19'b0000010_111101010110;
      15'b000_000111010101 : VALUE=19'b0000010_111101001001;
      15'b000_000111010110 : VALUE=19'b0000010_111100111100;
      15'b000_000111010111 : VALUE=19'b0000010_111100101111;
      15'b000_000111011000 : VALUE=19'b0000010_111100100010;
      15'b000_000111011001 : VALUE=19'b0000010_111100010101;
      15'b000_000111011010 : VALUE=19'b0000010_111100001001;
      15'b000_000111011011 : VALUE=19'b0000010_111011111100;
      15'b000_000111011100 : VALUE=19'b0000010_111011101111;
      15'b000_000111011101 : VALUE=19'b0000010_111011100011;
      15'b000_000111011110 : VALUE=19'b0000010_111011010110;
      15'b000_000111011111 : VALUE=19'b0000010_111011001010;
      15'b000_000111100000 : VALUE=19'b0000010_111010111101;
      15'b000_000111100001 : VALUE=19'b0000010_111010110001;
      15'b000_000111100010 : VALUE=19'b0000010_111010100100;
      15'b000_000111100011 : VALUE=19'b0000010_111010011000;
      15'b000_000111100100 : VALUE=19'b0000010_111010001100;
      15'b000_000111100101 : VALUE=19'b0000010_111001111111;
      15'b000_000111100110 : VALUE=19'b0000010_111001110011;
      15'b000_000111100111 : VALUE=19'b0000010_111001100111;
      15'b000_000111101000 : VALUE=19'b0000010_111001011011;
      15'b000_000111101001 : VALUE=19'b0000010_111001001111;
      15'b000_000111101010 : VALUE=19'b0000010_111001000010;
      15'b000_000111101011 : VALUE=19'b0000010_111000110110;
      15'b000_000111101100 : VALUE=19'b0000010_111000101010;
      15'b000_000111101101 : VALUE=19'b0000010_111000011110;
      15'b000_000111101110 : VALUE=19'b0000010_111000010010;
      15'b000_000111101111 : VALUE=19'b0000010_111000000110;
      15'b000_000111110000 : VALUE=19'b0000010_110111111011;
      15'b000_000111110001 : VALUE=19'b0000010_110111101111;
      15'b000_000111110010 : VALUE=19'b0000010_110111100011;
      15'b000_000111110011 : VALUE=19'b0000010_110111010111;
      15'b000_000111110100 : VALUE=19'b0000010_110111001011;
      15'b000_000111110101 : VALUE=19'b0000010_110111000000;
      15'b000_000111110110 : VALUE=19'b0000010_110110110100;
      15'b000_000111110111 : VALUE=19'b0000010_110110101000;
      15'b000_000111111000 : VALUE=19'b0000010_110110011101;
      15'b000_000111111001 : VALUE=19'b0000010_110110010001;
      15'b000_000111111010 : VALUE=19'b0000010_110110000110;
      15'b000_000111111011 : VALUE=19'b0000010_110101111010;
      15'b000_000111111100 : VALUE=19'b0000010_110101101111;
      15'b000_000111111101 : VALUE=19'b0000010_110101100011;
      15'b000_000111111110 : VALUE=19'b0000010_110101011000;
      15'b000_000111111111 : VALUE=19'b0000010_110101001101;
      15'b000_001000000000 : VALUE=19'b0000010_110101000001;
      15'b000_001000000001 : VALUE=19'b0000010_110100110110;
      15'b000_001000000010 : VALUE=19'b0000010_110100101011;
      15'b000_001000000011 : VALUE=19'b0000010_110100011111;
      15'b000_001000000100 : VALUE=19'b0000010_110100010100;
      15'b000_001000000101 : VALUE=19'b0000010_110100001001;
      15'b000_001000000110 : VALUE=19'b0000010_110011111110;
      15'b000_001000000111 : VALUE=19'b0000010_110011110011;
      15'b000_001000001000 : VALUE=19'b0000010_110011101000;
      15'b000_001000001001 : VALUE=19'b0000010_110011011101;
      15'b000_001000001010 : VALUE=19'b0000010_110011010010;
      15'b000_001000001011 : VALUE=19'b0000010_110011000111;
      15'b000_001000001100 : VALUE=19'b0000010_110010111100;
      15'b000_001000001101 : VALUE=19'b0000010_110010110001;
      15'b000_001000001110 : VALUE=19'b0000010_110010100110;
      15'b000_001000001111 : VALUE=19'b0000010_110010011011;
      15'b000_001000010000 : VALUE=19'b0000010_110010010000;
      15'b000_001000010001 : VALUE=19'b0000010_110010000110;
      15'b000_001000010010 : VALUE=19'b0000010_110001111011;
      15'b000_001000010011 : VALUE=19'b0000010_110001110000;
      15'b000_001000010100 : VALUE=19'b0000010_110001100101;
      15'b000_001000010101 : VALUE=19'b0000010_110001011011;
      15'b000_001000010110 : VALUE=19'b0000010_110001010000;
      15'b000_001000010111 : VALUE=19'b0000010_110001000101;
      15'b000_001000011000 : VALUE=19'b0000010_110000111011;
      15'b000_001000011001 : VALUE=19'b0000010_110000110000;
      15'b000_001000011010 : VALUE=19'b0000010_110000100110;
      15'b000_001000011011 : VALUE=19'b0000010_110000011011;
      15'b000_001000011100 : VALUE=19'b0000010_110000010001;
      15'b000_001000011101 : VALUE=19'b0000010_110000000110;
      15'b000_001000011110 : VALUE=19'b0000010_101111111100;
      15'b000_001000011111 : VALUE=19'b0000010_101111110010;
      15'b000_001000100000 : VALUE=19'b0000010_101111100111;
      15'b000_001000100001 : VALUE=19'b0000010_101111011101;
      15'b000_001000100010 : VALUE=19'b0000010_101111010011;
      15'b000_001000100011 : VALUE=19'b0000010_101111001000;
      15'b000_001000100100 : VALUE=19'b0000010_101110111110;
      15'b000_001000100101 : VALUE=19'b0000010_101110110100;
      15'b000_001000100110 : VALUE=19'b0000010_101110101010;
      15'b000_001000100111 : VALUE=19'b0000010_101110100000;
      15'b000_001000101000 : VALUE=19'b0000010_101110010110;
      15'b000_001000101001 : VALUE=19'b0000010_101110001011;
      15'b000_001000101010 : VALUE=19'b0000010_101110000001;
      15'b000_001000101011 : VALUE=19'b0000010_101101110111;
      15'b000_001000101100 : VALUE=19'b0000010_101101101101;
      15'b000_001000101101 : VALUE=19'b0000010_101101100011;
      15'b000_001000101110 : VALUE=19'b0000010_101101011001;
      15'b000_001000101111 : VALUE=19'b0000010_101101010000;
      15'b000_001000110000 : VALUE=19'b0000010_101101000110;
      15'b000_001000110001 : VALUE=19'b0000010_101100111100;
      15'b000_001000110010 : VALUE=19'b0000010_101100110010;
      15'b000_001000110011 : VALUE=19'b0000010_101100101000;
      15'b000_001000110100 : VALUE=19'b0000010_101100011110;
      15'b000_001000110101 : VALUE=19'b0000010_101100010100;
      15'b000_001000110110 : VALUE=19'b0000010_101100001011;
      15'b000_001000110111 : VALUE=19'b0000010_101100000001;
      15'b000_001000111000 : VALUE=19'b0000010_101011110111;
      15'b000_001000111001 : VALUE=19'b0000010_101011101110;
      15'b000_001000111010 : VALUE=19'b0000010_101011100100;
      15'b000_001000111011 : VALUE=19'b0000010_101011011010;
      15'b000_001000111100 : VALUE=19'b0000010_101011010001;
      15'b000_001000111101 : VALUE=19'b0000010_101011000111;
      15'b000_001000111110 : VALUE=19'b0000010_101010111110;
      15'b000_001000111111 : VALUE=19'b0000010_101010110100;
      15'b000_001001000000 : VALUE=19'b0000010_101010101011;
      15'b000_001001000001 : VALUE=19'b0000010_101010100001;
      15'b000_001001000010 : VALUE=19'b0000010_101010011000;
      15'b000_001001000011 : VALUE=19'b0000010_101010001110;
      15'b000_001001000100 : VALUE=19'b0000010_101010000101;
      15'b000_001001000101 : VALUE=19'b0000010_101001111100;
      15'b000_001001000110 : VALUE=19'b0000010_101001110010;
      15'b000_001001000111 : VALUE=19'b0000010_101001101001;
      15'b000_001001001000 : VALUE=19'b0000010_101001100000;
      15'b000_001001001001 : VALUE=19'b0000010_101001010110;
      15'b000_001001001010 : VALUE=19'b0000010_101001001101;
      15'b000_001001001011 : VALUE=19'b0000010_101001000100;
      15'b000_001001001100 : VALUE=19'b0000010_101000111011;
      15'b000_001001001101 : VALUE=19'b0000010_101000110001;
      15'b000_001001001110 : VALUE=19'b0000010_101000101000;
      15'b000_001001001111 : VALUE=19'b0000010_101000011111;
      15'b000_001001010000 : VALUE=19'b0000010_101000010110;
      15'b000_001001010001 : VALUE=19'b0000010_101000001101;
      15'b000_001001010010 : VALUE=19'b0000010_101000000100;
      15'b000_001001010011 : VALUE=19'b0000010_100111111011;
      15'b000_001001010100 : VALUE=19'b0000010_100111110010;
      15'b000_001001010101 : VALUE=19'b0000010_100111101001;
      15'b000_001001010110 : VALUE=19'b0000010_100111100000;
      15'b000_001001010111 : VALUE=19'b0000010_100111010111;
      15'b000_001001011000 : VALUE=19'b0000010_100111001110;
      15'b000_001001011001 : VALUE=19'b0000010_100111000101;
      15'b000_001001011010 : VALUE=19'b0000010_100110111100;
      15'b000_001001011011 : VALUE=19'b0000010_100110110011;
      15'b000_001001011100 : VALUE=19'b0000010_100110101010;
      15'b000_001001011101 : VALUE=19'b0000010_100110100010;
      15'b000_001001011110 : VALUE=19'b0000010_100110011001;
      15'b000_001001011111 : VALUE=19'b0000010_100110010000;
      15'b000_001001100000 : VALUE=19'b0000010_100110000111;
      15'b000_001001100001 : VALUE=19'b0000010_100101111111;
      15'b000_001001100010 : VALUE=19'b0000010_100101110110;
      15'b000_001001100011 : VALUE=19'b0000010_100101101101;
      15'b000_001001100100 : VALUE=19'b0000010_100101100101;
      15'b000_001001100101 : VALUE=19'b0000010_100101011100;
      15'b000_001001100110 : VALUE=19'b0000010_100101010011;
      15'b000_001001100111 : VALUE=19'b0000010_100101001011;
      15'b000_001001101000 : VALUE=19'b0000010_100101000010;
      15'b000_001001101001 : VALUE=19'b0000010_100100111010;
      15'b000_001001101010 : VALUE=19'b0000010_100100110001;
      15'b000_001001101011 : VALUE=19'b0000010_100100101000;
      15'b000_001001101100 : VALUE=19'b0000010_100100100000;
      15'b000_001001101101 : VALUE=19'b0000010_100100010111;
      15'b000_001001101110 : VALUE=19'b0000010_100100001111;
      15'b000_001001101111 : VALUE=19'b0000010_100100000111;
      15'b000_001001110000 : VALUE=19'b0000010_100011111110;
      15'b000_001001110001 : VALUE=19'b0000010_100011110110;
      15'b000_001001110010 : VALUE=19'b0000010_100011101101;
      15'b000_001001110011 : VALUE=19'b0000010_100011100101;
      15'b000_001001110100 : VALUE=19'b0000010_100011011101;
      15'b000_001001110101 : VALUE=19'b0000010_100011010100;
      15'b000_001001110110 : VALUE=19'b0000010_100011001100;
      15'b000_001001110111 : VALUE=19'b0000010_100011000100;
      15'b000_001001111000 : VALUE=19'b0000010_100010111100;
      15'b000_001001111001 : VALUE=19'b0000010_100010110011;
      15'b000_001001111010 : VALUE=19'b0000010_100010101011;
      15'b000_001001111011 : VALUE=19'b0000010_100010100011;
      15'b000_001001111100 : VALUE=19'b0000010_100010011011;
      15'b000_001001111101 : VALUE=19'b0000010_100010010011;
      15'b000_001001111110 : VALUE=19'b0000010_100010001010;
      15'b000_001001111111 : VALUE=19'b0000010_100010000010;
      15'b000_001010000000 : VALUE=19'b0000010_100001111010;
      15'b000_001010000001 : VALUE=19'b0000010_100001110010;
      15'b000_001010000010 : VALUE=19'b0000010_100001101010;
      15'b000_001010000011 : VALUE=19'b0000010_100001100010;
      15'b000_001010000100 : VALUE=19'b0000010_100001011010;
      15'b000_001010000101 : VALUE=19'b0000010_100001010010;
      15'b000_001010000110 : VALUE=19'b0000010_100001001010;
      15'b000_001010000111 : VALUE=19'b0000010_100001000010;
      15'b000_001010001000 : VALUE=19'b0000010_100000111010;
      15'b000_001010001001 : VALUE=19'b0000010_100000110010;
      15'b000_001010001010 : VALUE=19'b0000010_100000101010;
      15'b000_001010001011 : VALUE=19'b0000010_100000100010;
      15'b000_001010001100 : VALUE=19'b0000010_100000011010;
      15'b000_001010001101 : VALUE=19'b0000010_100000010010;
      15'b000_001010001110 : VALUE=19'b0000010_100000001011;
      15'b000_001010001111 : VALUE=19'b0000010_100000000011;
      15'b000_001010010000 : VALUE=19'b0000010_011111111011;
      15'b000_001010010001 : VALUE=19'b0000010_011111110011;
      15'b000_001010010010 : VALUE=19'b0000010_011111101011;
      15'b000_001010010011 : VALUE=19'b0000010_011111100100;
      15'b000_001010010100 : VALUE=19'b0000010_011111011100;
      15'b000_001010010101 : VALUE=19'b0000010_011111010100;
      15'b000_001010010110 : VALUE=19'b0000010_011111001101;
      15'b000_001010010111 : VALUE=19'b0000010_011111000101;
      15'b000_001010011000 : VALUE=19'b0000010_011110111101;
      15'b000_001010011001 : VALUE=19'b0000010_011110110110;
      15'b000_001010011010 : VALUE=19'b0000010_011110101110;
      15'b000_001010011011 : VALUE=19'b0000010_011110100110;
      15'b000_001010011100 : VALUE=19'b0000010_011110011111;
      15'b000_001010011101 : VALUE=19'b0000010_011110010111;
      15'b000_001010011110 : VALUE=19'b0000010_011110010000;
      15'b000_001010011111 : VALUE=19'b0000010_011110001000;
      15'b000_001010100000 : VALUE=19'b0000010_011110000000;
      15'b000_001010100001 : VALUE=19'b0000010_011101111001;
      15'b000_001010100010 : VALUE=19'b0000010_011101110001;
      15'b000_001010100011 : VALUE=19'b0000010_011101101010;
      15'b000_001010100100 : VALUE=19'b0000010_011101100010;
      15'b000_001010100101 : VALUE=19'b0000010_011101011011;
      15'b000_001010100110 : VALUE=19'b0000010_011101010100;
      15'b000_001010100111 : VALUE=19'b0000010_011101001100;
      15'b000_001010101000 : VALUE=19'b0000010_011101000101;
      15'b000_001010101001 : VALUE=19'b0000010_011100111101;
      15'b000_001010101010 : VALUE=19'b0000010_011100110110;
      15'b000_001010101011 : VALUE=19'b0000010_011100101111;
      15'b000_001010101100 : VALUE=19'b0000010_011100100111;
      15'b000_001010101101 : VALUE=19'b0000010_011100100000;
      15'b000_001010101110 : VALUE=19'b0000010_011100011001;
      15'b000_001010101111 : VALUE=19'b0000010_011100010001;
      15'b000_001010110000 : VALUE=19'b0000010_011100001010;
      15'b000_001010110001 : VALUE=19'b0000010_011100000011;
      15'b000_001010110010 : VALUE=19'b0000010_011011111100;
      15'b000_001010110011 : VALUE=19'b0000010_011011110100;
      15'b000_001010110100 : VALUE=19'b0000010_011011101101;
      15'b000_001010110101 : VALUE=19'b0000010_011011100110;
      15'b000_001010110110 : VALUE=19'b0000010_011011011111;
      15'b000_001010110111 : VALUE=19'b0000010_011011011000;
      15'b000_001010111000 : VALUE=19'b0000010_011011010001;
      15'b000_001010111001 : VALUE=19'b0000010_011011001001;
      15'b000_001010111010 : VALUE=19'b0000010_011011000010;
      15'b000_001010111011 : VALUE=19'b0000010_011010111011;
      15'b000_001010111100 : VALUE=19'b0000010_011010110100;
      15'b000_001010111101 : VALUE=19'b0000010_011010101101;
      15'b000_001010111110 : VALUE=19'b0000010_011010100110;
      15'b000_001010111111 : VALUE=19'b0000010_011010011111;
      15'b000_001011000000 : VALUE=19'b0000010_011010011000;
      15'b000_001011000001 : VALUE=19'b0000010_011010010001;
      15'b000_001011000010 : VALUE=19'b0000010_011010001010;
      15'b000_001011000011 : VALUE=19'b0000010_011010000011;
      15'b000_001011000100 : VALUE=19'b0000010_011001111100;
      15'b000_001011000101 : VALUE=19'b0000010_011001110101;
      15'b000_001011000110 : VALUE=19'b0000010_011001101110;
      15'b000_001011000111 : VALUE=19'b0000010_011001100111;
      15'b000_001011001000 : VALUE=19'b0000010_011001100000;
      15'b000_001011001001 : VALUE=19'b0000010_011001011001;
      15'b000_001011001010 : VALUE=19'b0000010_011001010010;
      15'b000_001011001011 : VALUE=19'b0000010_011001001100;
      15'b000_001011001100 : VALUE=19'b0000010_011001000101;
      15'b000_001011001101 : VALUE=19'b0000010_011000111110;
      15'b000_001011001110 : VALUE=19'b0000010_011000110111;
      15'b000_001011001111 : VALUE=19'b0000010_011000110000;
      15'b000_001011010000 : VALUE=19'b0000010_011000101010;
      15'b000_001011010001 : VALUE=19'b0000010_011000100011;
      15'b000_001011010010 : VALUE=19'b0000010_011000011100;
      15'b000_001011010011 : VALUE=19'b0000010_011000010101;
      15'b000_001011010100 : VALUE=19'b0000010_011000001111;
      15'b000_001011010101 : VALUE=19'b0000010_011000001000;
      15'b000_001011010110 : VALUE=19'b0000010_011000000001;
      15'b000_001011010111 : VALUE=19'b0000010_010111111010;
      15'b000_001011011000 : VALUE=19'b0000010_010111110100;
      15'b000_001011011001 : VALUE=19'b0000010_010111101101;
      15'b000_001011011010 : VALUE=19'b0000010_010111100110;
      15'b000_001011011011 : VALUE=19'b0000010_010111100000;
      15'b000_001011011100 : VALUE=19'b0000010_010111011001;
      15'b000_001011011101 : VALUE=19'b0000010_010111010011;
      15'b000_001011011110 : VALUE=19'b0000010_010111001100;
      15'b000_001011011111 : VALUE=19'b0000010_010111000101;
      15'b000_001011100000 : VALUE=19'b0000010_010110111111;
      15'b000_001011100001 : VALUE=19'b0000010_010110111000;
      15'b000_001011100010 : VALUE=19'b0000010_010110110010;
      15'b000_001011100011 : VALUE=19'b0000010_010110101011;
      15'b000_001011100100 : VALUE=19'b0000010_010110100101;
      15'b000_001011100101 : VALUE=19'b0000010_010110011110;
      15'b000_001011100110 : VALUE=19'b0000010_010110011000;
      15'b000_001011100111 : VALUE=19'b0000010_010110010001;
      15'b000_001011101000 : VALUE=19'b0000010_010110001011;
      15'b000_001011101001 : VALUE=19'b0000010_010110000100;
      15'b000_001011101010 : VALUE=19'b0000010_010101111110;
      15'b000_001011101011 : VALUE=19'b0000010_010101110111;
      15'b000_001011101100 : VALUE=19'b0000010_010101110001;
      15'b000_001011101101 : VALUE=19'b0000010_010101101011;
      15'b000_001011101110 : VALUE=19'b0000010_010101100100;
      15'b000_001011101111 : VALUE=19'b0000010_010101011110;
      15'b000_001011110000 : VALUE=19'b0000010_010101010111;
      15'b000_001011110001 : VALUE=19'b0000010_010101010001;
      15'b000_001011110010 : VALUE=19'b0000010_010101001011;
      15'b000_001011110011 : VALUE=19'b0000010_010101000100;
      15'b000_001011110100 : VALUE=19'b0000010_010100111110;
      15'b000_001011110101 : VALUE=19'b0000010_010100111000;
      15'b000_001011110110 : VALUE=19'b0000010_010100110001;
      15'b000_001011110111 : VALUE=19'b0000010_010100101011;
      15'b000_001011111000 : VALUE=19'b0000010_010100100101;
      15'b000_001011111001 : VALUE=19'b0000010_010100011111;
      15'b000_001011111010 : VALUE=19'b0000010_010100011000;
      15'b000_001011111011 : VALUE=19'b0000010_010100010010;
      15'b000_001011111100 : VALUE=19'b0000010_010100001100;
      15'b000_001011111101 : VALUE=19'b0000010_010100000110;
      15'b000_001011111110 : VALUE=19'b0000010_010100000000;
      15'b000_001011111111 : VALUE=19'b0000010_010011111001;
      15'b000_001100000000 : VALUE=19'b0000010_010011110011;
      15'b000_001100000001 : VALUE=19'b0000010_010011101101;
      15'b000_001100000010 : VALUE=19'b0000010_010011100111;
      15'b000_001100000011 : VALUE=19'b0000010_010011100001;
      15'b000_001100000100 : VALUE=19'b0000010_010011011011;
      15'b000_001100000101 : VALUE=19'b0000010_010011010101;
      15'b000_001100000110 : VALUE=19'b0000010_010011001111;
      15'b000_001100000111 : VALUE=19'b0000010_010011001000;
      15'b000_001100001000 : VALUE=19'b0000010_010011000010;
      15'b000_001100001001 : VALUE=19'b0000010_010010111100;
      15'b000_001100001010 : VALUE=19'b0000010_010010110110;
      15'b000_001100001011 : VALUE=19'b0000010_010010110000;
      15'b000_001100001100 : VALUE=19'b0000010_010010101010;
      15'b000_001100001101 : VALUE=19'b0000010_010010100100;
      15'b000_001100001110 : VALUE=19'b0000010_010010011110;
      15'b000_001100001111 : VALUE=19'b0000010_010010011000;
      15'b000_001100010000 : VALUE=19'b0000010_010010010010;
      15'b000_001100010001 : VALUE=19'b0000010_010010001100;
      15'b000_001100010010 : VALUE=19'b0000010_010010000110;
      15'b000_001100010011 : VALUE=19'b0000010_010010000000;
      15'b000_001100010100 : VALUE=19'b0000010_010001111010;
      15'b000_001100010101 : VALUE=19'b0000010_010001110101;
      15'b000_001100010110 : VALUE=19'b0000010_010001101111;
      15'b000_001100010111 : VALUE=19'b0000010_010001101001;
      15'b000_001100011000 : VALUE=19'b0000010_010001100011;
      15'b000_001100011001 : VALUE=19'b0000010_010001011101;
      15'b000_001100011010 : VALUE=19'b0000010_010001010111;
      15'b000_001100011011 : VALUE=19'b0000010_010001010001;
      15'b000_001100011100 : VALUE=19'b0000010_010001001011;
      15'b000_001100011101 : VALUE=19'b0000010_010001000110;
      15'b000_001100011110 : VALUE=19'b0000010_010001000000;
      15'b000_001100011111 : VALUE=19'b0000010_010000111010;
      15'b000_001100100000 : VALUE=19'b0000010_010000110100;
      15'b000_001100100001 : VALUE=19'b0000010_010000101110;
      15'b000_001100100010 : VALUE=19'b0000010_010000101001;
      15'b000_001100100011 : VALUE=19'b0000010_010000100011;
      15'b000_001100100100 : VALUE=19'b0000010_010000011101;
      15'b000_001100100101 : VALUE=19'b0000010_010000010111;
      15'b000_001100100110 : VALUE=19'b0000010_010000010010;
      15'b000_001100100111 : VALUE=19'b0000010_010000001100;
      15'b000_001100101000 : VALUE=19'b0000010_010000000110;
      15'b000_001100101001 : VALUE=19'b0000010_010000000000;
      15'b000_001100101010 : VALUE=19'b0000010_001111111011;
      15'b000_001100101011 : VALUE=19'b0000010_001111110101;
      15'b000_001100101100 : VALUE=19'b0000010_001111101111;
      15'b000_001100101101 : VALUE=19'b0000010_001111101010;
      15'b000_001100101110 : VALUE=19'b0000010_001111100100;
      15'b000_001100101111 : VALUE=19'b0000010_001111011111;
      15'b000_001100110000 : VALUE=19'b0000010_001111011001;
      15'b000_001100110001 : VALUE=19'b0000010_001111010011;
      15'b000_001100110010 : VALUE=19'b0000010_001111001110;
      15'b000_001100110011 : VALUE=19'b0000010_001111001000;
      15'b000_001100110100 : VALUE=19'b0000010_001111000010;
      15'b000_001100110101 : VALUE=19'b0000010_001110111101;
      15'b000_001100110110 : VALUE=19'b0000010_001110110111;
      15'b000_001100110111 : VALUE=19'b0000010_001110110010;
      15'b000_001100111000 : VALUE=19'b0000010_001110101100;
      15'b000_001100111001 : VALUE=19'b0000010_001110100111;
      15'b000_001100111010 : VALUE=19'b0000010_001110100001;
      15'b000_001100111011 : VALUE=19'b0000010_001110011100;
      15'b000_001100111100 : VALUE=19'b0000010_001110010110;
      15'b000_001100111101 : VALUE=19'b0000010_001110010001;
      15'b000_001100111110 : VALUE=19'b0000010_001110001011;
      15'b000_001100111111 : VALUE=19'b0000010_001110000110;
      15'b000_001101000000 : VALUE=19'b0000010_001110000000;
      15'b000_001101000001 : VALUE=19'b0000010_001101111011;
      15'b000_001101000010 : VALUE=19'b0000010_001101110101;
      15'b000_001101000011 : VALUE=19'b0000010_001101110000;
      15'b000_001101000100 : VALUE=19'b0000010_001101101010;
      15'b000_001101000101 : VALUE=19'b0000010_001101100101;
      15'b000_001101000110 : VALUE=19'b0000010_001101100000;
      15'b000_001101000111 : VALUE=19'b0000010_001101011010;
      15'b000_001101001000 : VALUE=19'b0000010_001101010101;
      15'b000_001101001001 : VALUE=19'b0000010_001101001111;
      15'b000_001101001010 : VALUE=19'b0000010_001101001010;
      15'b000_001101001011 : VALUE=19'b0000010_001101000101;
      15'b000_001101001100 : VALUE=19'b0000010_001100111111;
      15'b000_001101001101 : VALUE=19'b0000010_001100111010;
      15'b000_001101001110 : VALUE=19'b0000010_001100110101;
      15'b000_001101001111 : VALUE=19'b0000010_001100101111;
      15'b000_001101010000 : VALUE=19'b0000010_001100101010;
      15'b000_001101010001 : VALUE=19'b0000010_001100100101;
      15'b000_001101010010 : VALUE=19'b0000010_001100011111;
      15'b000_001101010011 : VALUE=19'b0000010_001100011010;
      15'b000_001101010100 : VALUE=19'b0000010_001100010101;
      15'b000_001101010101 : VALUE=19'b0000010_001100010000;
      15'b000_001101010110 : VALUE=19'b0000010_001100001010;
      15'b000_001101010111 : VALUE=19'b0000010_001100000101;
      15'b000_001101011000 : VALUE=19'b0000010_001100000000;
      15'b000_001101011001 : VALUE=19'b0000010_001011111011;
      15'b000_001101011010 : VALUE=19'b0000010_001011110101;
      15'b000_001101011011 : VALUE=19'b0000010_001011110000;
      15'b000_001101011100 : VALUE=19'b0000010_001011101011;
      15'b000_001101011101 : VALUE=19'b0000010_001011100110;
      15'b000_001101011110 : VALUE=19'b0000010_001011100001;
      15'b000_001101011111 : VALUE=19'b0000010_001011011011;
      15'b000_001101100000 : VALUE=19'b0000010_001011010110;
      15'b000_001101100001 : VALUE=19'b0000010_001011010001;
      15'b000_001101100010 : VALUE=19'b0000010_001011001100;
      15'b000_001101100011 : VALUE=19'b0000010_001011000111;
      15'b000_001101100100 : VALUE=19'b0000010_001011000010;
      15'b000_001101100101 : VALUE=19'b0000010_001010111101;
      15'b000_001101100110 : VALUE=19'b0000010_001010111000;
      15'b000_001101100111 : VALUE=19'b0000010_001010110010;
      15'b000_001101101000 : VALUE=19'b0000010_001010101101;
      15'b000_001101101001 : VALUE=19'b0000010_001010101000;
      15'b000_001101101010 : VALUE=19'b0000010_001010100011;
      15'b000_001101101011 : VALUE=19'b0000010_001010011110;
      15'b000_001101101100 : VALUE=19'b0000010_001010011001;
      15'b000_001101101101 : VALUE=19'b0000010_001010010100;
      15'b000_001101101110 : VALUE=19'b0000010_001010001111;
      15'b000_001101101111 : VALUE=19'b0000010_001010001010;
      15'b000_001101110000 : VALUE=19'b0000010_001010000101;
      15'b000_001101110001 : VALUE=19'b0000010_001010000000;
      15'b000_001101110010 : VALUE=19'b0000010_001001111011;
      15'b000_001101110011 : VALUE=19'b0000010_001001110110;
      15'b000_001101110100 : VALUE=19'b0000010_001001110001;
      15'b000_001101110101 : VALUE=19'b0000010_001001101100;
      15'b000_001101110110 : VALUE=19'b0000010_001001100111;
      15'b000_001101110111 : VALUE=19'b0000010_001001100010;
      15'b000_001101111000 : VALUE=19'b0000010_001001011101;
      15'b000_001101111001 : VALUE=19'b0000010_001001011000;
      15'b000_001101111010 : VALUE=19'b0000010_001001010011;
      15'b000_001101111011 : VALUE=19'b0000010_001001001110;
      15'b000_001101111100 : VALUE=19'b0000010_001001001001;
      15'b000_001101111101 : VALUE=19'b0000010_001001000100;
      15'b000_001101111110 : VALUE=19'b0000010_001000111111;
      15'b000_001101111111 : VALUE=19'b0000010_001000111011;
      15'b000_001110000000 : VALUE=19'b0000010_001000110110;
      15'b000_001110000001 : VALUE=19'b0000010_001000110001;
      15'b000_001110000010 : VALUE=19'b0000010_001000101100;
      15'b000_001110000011 : VALUE=19'b0000010_001000100111;
      15'b000_001110000100 : VALUE=19'b0000010_001000100010;
      15'b000_001110000101 : VALUE=19'b0000010_001000011101;
      15'b000_001110000110 : VALUE=19'b0000010_001000011000;
      15'b000_001110000111 : VALUE=19'b0000010_001000010100;
      15'b000_001110001000 : VALUE=19'b0000010_001000001111;
      15'b000_001110001001 : VALUE=19'b0000010_001000001010;
      15'b000_001110001010 : VALUE=19'b0000010_001000000101;
      15'b000_001110001011 : VALUE=19'b0000010_001000000000;
      15'b000_001110001100 : VALUE=19'b0000010_000111111100;
      15'b000_001110001101 : VALUE=19'b0000010_000111110111;
      15'b000_001110001110 : VALUE=19'b0000010_000111110010;
      15'b000_001110001111 : VALUE=19'b0000010_000111101101;
      15'b000_001110010000 : VALUE=19'b0000010_000111101000;
      15'b000_001110010001 : VALUE=19'b0000010_000111100100;
      15'b000_001110010010 : VALUE=19'b0000010_000111011111;
      15'b000_001110010011 : VALUE=19'b0000010_000111011010;
      15'b000_001110010100 : VALUE=19'b0000010_000111010101;
      15'b000_001110010101 : VALUE=19'b0000010_000111010001;
      15'b000_001110010110 : VALUE=19'b0000010_000111001100;
      15'b000_001110010111 : VALUE=19'b0000010_000111000111;
      15'b000_001110011000 : VALUE=19'b0000010_000111000011;
      15'b000_001110011001 : VALUE=19'b0000010_000110111110;
      15'b000_001110011010 : VALUE=19'b0000010_000110111001;
      15'b000_001110011011 : VALUE=19'b0000010_000110110101;
      15'b000_001110011100 : VALUE=19'b0000010_000110110000;
      15'b000_001110011101 : VALUE=19'b0000010_000110101011;
      15'b000_001110011110 : VALUE=19'b0000010_000110100111;
      15'b000_001110011111 : VALUE=19'b0000010_000110100010;
      15'b000_001110100000 : VALUE=19'b0000010_000110011101;
      15'b000_001110100001 : VALUE=19'b0000010_000110011001;
      15'b000_001110100010 : VALUE=19'b0000010_000110010100;
      15'b000_001110100011 : VALUE=19'b0000010_000110001111;
      15'b000_001110100100 : VALUE=19'b0000010_000110001011;
      15'b000_001110100101 : VALUE=19'b0000010_000110000110;
      15'b000_001110100110 : VALUE=19'b0000010_000110000010;
      15'b000_001110100111 : VALUE=19'b0000010_000101111101;
      15'b000_001110101000 : VALUE=19'b0000010_000101111000;
      15'b000_001110101001 : VALUE=19'b0000010_000101110100;
      15'b000_001110101010 : VALUE=19'b0000010_000101101111;
      15'b000_001110101011 : VALUE=19'b0000010_000101101011;
      15'b000_001110101100 : VALUE=19'b0000010_000101100110;
      15'b000_001110101101 : VALUE=19'b0000010_000101100010;
      15'b000_001110101110 : VALUE=19'b0000010_000101011101;
      15'b000_001110101111 : VALUE=19'b0000010_000101011001;
      15'b000_001110110000 : VALUE=19'b0000010_000101010100;
      15'b000_001110110001 : VALUE=19'b0000010_000101010000;
      15'b000_001110110010 : VALUE=19'b0000010_000101001011;
      15'b000_001110110011 : VALUE=19'b0000010_000101000111;
      15'b000_001110110100 : VALUE=19'b0000010_000101000010;
      15'b000_001110110101 : VALUE=19'b0000010_000100111110;
      15'b000_001110110110 : VALUE=19'b0000010_000100111001;
      15'b000_001110110111 : VALUE=19'b0000010_000100110101;
      15'b000_001110111000 : VALUE=19'b0000010_000100110000;
      15'b000_001110111001 : VALUE=19'b0000010_000100101100;
      15'b000_001110111010 : VALUE=19'b0000010_000100100111;
      15'b000_001110111011 : VALUE=19'b0000010_000100100011;
      15'b000_001110111100 : VALUE=19'b0000010_000100011110;
      15'b000_001110111101 : VALUE=19'b0000010_000100011010;
      15'b000_001110111110 : VALUE=19'b0000010_000100010101;
      15'b000_001110111111 : VALUE=19'b0000010_000100010001;
      15'b000_001111000000 : VALUE=19'b0000010_000100001101;
      15'b000_001111000001 : VALUE=19'b0000010_000100001000;
      15'b000_001111000010 : VALUE=19'b0000010_000100000100;
      15'b000_001111000011 : VALUE=19'b0000010_000011111111;
      15'b000_001111000100 : VALUE=19'b0000010_000011111011;
      15'b000_001111000101 : VALUE=19'b0000010_000011110111;
      15'b000_001111000110 : VALUE=19'b0000010_000011110010;
      15'b000_001111000111 : VALUE=19'b0000010_000011101110;
      15'b000_001111001000 : VALUE=19'b0000010_000011101010;
      15'b000_001111001001 : VALUE=19'b0000010_000011100101;
      15'b000_001111001010 : VALUE=19'b0000010_000011100001;
      15'b000_001111001011 : VALUE=19'b0000010_000011011101;
      15'b000_001111001100 : VALUE=19'b0000010_000011011000;
      15'b000_001111001101 : VALUE=19'b0000010_000011010100;
      15'b000_001111001110 : VALUE=19'b0000010_000011010000;
      15'b000_001111001111 : VALUE=19'b0000010_000011001011;
      15'b000_001111010000 : VALUE=19'b0000010_000011000111;
      15'b000_001111010001 : VALUE=19'b0000010_000011000011;
      15'b000_001111010010 : VALUE=19'b0000010_000010111110;
      15'b000_001111010011 : VALUE=19'b0000010_000010111010;
      15'b000_001111010100 : VALUE=19'b0000010_000010110110;
      15'b000_001111010101 : VALUE=19'b0000010_000010110010;
      15'b000_001111010110 : VALUE=19'b0000010_000010101101;
      15'b000_001111010111 : VALUE=19'b0000010_000010101001;
      15'b000_001111011000 : VALUE=19'b0000010_000010100101;
      15'b000_001111011001 : VALUE=19'b0000010_000010100001;
      15'b000_001111011010 : VALUE=19'b0000010_000010011100;
      15'b000_001111011011 : VALUE=19'b0000010_000010011000;
      15'b000_001111011100 : VALUE=19'b0000010_000010010100;
      15'b000_001111011101 : VALUE=19'b0000010_000010010000;
      15'b000_001111011110 : VALUE=19'b0000010_000010001011;
      15'b000_001111011111 : VALUE=19'b0000010_000010000111;
      15'b000_001111100000 : VALUE=19'b0000010_000010000011;
      15'b000_001111100001 : VALUE=19'b0000010_000001111111;
      15'b000_001111100010 : VALUE=19'b0000010_000001111011;
      15'b000_001111100011 : VALUE=19'b0000010_000001110111;
      15'b000_001111100100 : VALUE=19'b0000010_000001110010;
      15'b000_001111100101 : VALUE=19'b0000010_000001101110;
      15'b000_001111100110 : VALUE=19'b0000010_000001101010;
      15'b000_001111100111 : VALUE=19'b0000010_000001100110;
      15'b000_001111101000 : VALUE=19'b0000010_000001100010;
      15'b000_001111101001 : VALUE=19'b0000010_000001011110;
      15'b000_001111101010 : VALUE=19'b0000010_000001011001;
      15'b000_001111101011 : VALUE=19'b0000010_000001010101;
      15'b000_001111101100 : VALUE=19'b0000010_000001010001;
      15'b000_001111101101 : VALUE=19'b0000010_000001001101;
      15'b000_001111101110 : VALUE=19'b0000010_000001001001;
      15'b000_001111101111 : VALUE=19'b0000010_000001000101;
      15'b000_001111110000 : VALUE=19'b0000010_000001000001;
      15'b000_001111110001 : VALUE=19'b0000010_000000111101;
      15'b000_001111110010 : VALUE=19'b0000010_000000111001;
      15'b000_001111110011 : VALUE=19'b0000010_000000110101;
      15'b000_001111110100 : VALUE=19'b0000010_000000110000;
      15'b000_001111110101 : VALUE=19'b0000010_000000101100;
      15'b000_001111110110 : VALUE=19'b0000010_000000101000;
      15'b000_001111110111 : VALUE=19'b0000010_000000100100;
      15'b000_001111111000 : VALUE=19'b0000010_000000100000;
      15'b000_001111111001 : VALUE=19'b0000010_000000011100;
      15'b000_001111111010 : VALUE=19'b0000010_000000011000;
      15'b000_001111111011 : VALUE=19'b0000010_000000010100;
      15'b000_001111111100 : VALUE=19'b0000010_000000010000;
      15'b000_001111111101 : VALUE=19'b0000010_000000001100;
      15'b000_001111111110 : VALUE=19'b0000010_000000001000;
      15'b000_001111111111 : VALUE=19'b0000010_000000000100;
      15'b000_010000000000 : VALUE=19'b0000010_000000000000;
      15'b000_010000000001 : VALUE=19'b0000001_111111111100;
      15'b000_010000000010 : VALUE=19'b0000001_111111111000;
      15'b000_010000000011 : VALUE=19'b0000001_111111110100;
      15'b000_010000000100 : VALUE=19'b0000001_111111110000;
      15'b000_010000000101 : VALUE=19'b0000001_111111101100;
      15'b000_010000000110 : VALUE=19'b0000001_111111101000;
      15'b000_010000000111 : VALUE=19'b0000001_111111100100;
      15'b000_010000001000 : VALUE=19'b0000001_111111100000;
      15'b000_010000001001 : VALUE=19'b0000001_111111011100;
      15'b000_010000001010 : VALUE=19'b0000001_111111011000;
      15'b000_010000001011 : VALUE=19'b0000001_111111010100;
      15'b000_010000001100 : VALUE=19'b0000001_111111010000;
      15'b000_010000001101 : VALUE=19'b0000001_111111001100;
      15'b000_010000001110 : VALUE=19'b0000001_111111001001;
      15'b000_010000001111 : VALUE=19'b0000001_111111000101;
      15'b000_010000010000 : VALUE=19'b0000001_111111000001;
      15'b000_010000010001 : VALUE=19'b0000001_111110111101;
      15'b000_010000010010 : VALUE=19'b0000001_111110111001;
      15'b000_010000010011 : VALUE=19'b0000001_111110110101;
      15'b000_010000010100 : VALUE=19'b0000001_111110110001;
      15'b000_010000010101 : VALUE=19'b0000001_111110101101;
      15'b000_010000010110 : VALUE=19'b0000001_111110101001;
      15'b000_010000010111 : VALUE=19'b0000001_111110100110;
      15'b000_010000011000 : VALUE=19'b0000001_111110100010;
      15'b000_010000011001 : VALUE=19'b0000001_111110011110;
      15'b000_010000011010 : VALUE=19'b0000001_111110011010;
      15'b000_010000011011 : VALUE=19'b0000001_111110010110;
      15'b000_010000011100 : VALUE=19'b0000001_111110010010;
      15'b000_010000011101 : VALUE=19'b0000001_111110001110;
      15'b000_010000011110 : VALUE=19'b0000001_111110001011;
      15'b000_010000011111 : VALUE=19'b0000001_111110000111;
      15'b000_010000100000 : VALUE=19'b0000001_111110000011;
      15'b000_010000100001 : VALUE=19'b0000001_111101111111;
      15'b000_010000100010 : VALUE=19'b0000001_111101111011;
      15'b000_010000100011 : VALUE=19'b0000001_111101110111;
      15'b000_010000100100 : VALUE=19'b0000001_111101110100;
      15'b000_010000100101 : VALUE=19'b0000001_111101110000;
      15'b000_010000100110 : VALUE=19'b0000001_111101101100;
      15'b000_010000100111 : VALUE=19'b0000001_111101101000;
      15'b000_010000101000 : VALUE=19'b0000001_111101100101;
      15'b000_010000101001 : VALUE=19'b0000001_111101100001;
      15'b000_010000101010 : VALUE=19'b0000001_111101011101;
      15'b000_010000101011 : VALUE=19'b0000001_111101011001;
      15'b000_010000101100 : VALUE=19'b0000001_111101010101;
      15'b000_010000101101 : VALUE=19'b0000001_111101010010;
      15'b000_010000101110 : VALUE=19'b0000001_111101001110;
      15'b000_010000101111 : VALUE=19'b0000001_111101001010;
      15'b000_010000110000 : VALUE=19'b0000001_111101000110;
      15'b000_010000110001 : VALUE=19'b0000001_111101000011;
      15'b000_010000110010 : VALUE=19'b0000001_111100111111;
      15'b000_010000110011 : VALUE=19'b0000001_111100111011;
      15'b000_010000110100 : VALUE=19'b0000001_111100111000;
      15'b000_010000110101 : VALUE=19'b0000001_111100110100;
      15'b000_010000110110 : VALUE=19'b0000001_111100110000;
      15'b000_010000110111 : VALUE=19'b0000001_111100101100;
      15'b000_010000111000 : VALUE=19'b0000001_111100101001;
      15'b000_010000111001 : VALUE=19'b0000001_111100100101;
      15'b000_010000111010 : VALUE=19'b0000001_111100100001;
      15'b000_010000111011 : VALUE=19'b0000001_111100011110;
      15'b000_010000111100 : VALUE=19'b0000001_111100011010;
      15'b000_010000111101 : VALUE=19'b0000001_111100010110;
      15'b000_010000111110 : VALUE=19'b0000001_111100010011;
      15'b000_010000111111 : VALUE=19'b0000001_111100001111;
      15'b000_010001000000 : VALUE=19'b0000001_111100001011;
      15'b000_010001000001 : VALUE=19'b0000001_111100001000;
      15'b000_010001000010 : VALUE=19'b0000001_111100000100;
      15'b000_010001000011 : VALUE=19'b0000001_111100000000;
      15'b000_010001000100 : VALUE=19'b0000001_111011111101;
      15'b000_010001000101 : VALUE=19'b0000001_111011111001;
      15'b000_010001000110 : VALUE=19'b0000001_111011110110;
      15'b000_010001000111 : VALUE=19'b0000001_111011110010;
      15'b000_010001001000 : VALUE=19'b0000001_111011101110;
      15'b000_010001001001 : VALUE=19'b0000001_111011101011;
      15'b000_010001001010 : VALUE=19'b0000001_111011100111;
      15'b000_010001001011 : VALUE=19'b0000001_111011100100;
      15'b000_010001001100 : VALUE=19'b0000001_111011100000;
      15'b000_010001001101 : VALUE=19'b0000001_111011011100;
      15'b000_010001001110 : VALUE=19'b0000001_111011011001;
      15'b000_010001001111 : VALUE=19'b0000001_111011010101;
      15'b000_010001010000 : VALUE=19'b0000001_111011010010;
      15'b000_010001010001 : VALUE=19'b0000001_111011001110;
      15'b000_010001010010 : VALUE=19'b0000001_111011001010;
      15'b000_010001010011 : VALUE=19'b0000001_111011000111;
      15'b000_010001010100 : VALUE=19'b0000001_111011000011;
      15'b000_010001010101 : VALUE=19'b0000001_111011000000;
      15'b000_010001010110 : VALUE=19'b0000001_111010111100;
      15'b000_010001010111 : VALUE=19'b0000001_111010111001;
      15'b000_010001011000 : VALUE=19'b0000001_111010110101;
      15'b000_010001011001 : VALUE=19'b0000001_111010110010;
      15'b000_010001011010 : VALUE=19'b0000001_111010101110;
      15'b000_010001011011 : VALUE=19'b0000001_111010101011;
      15'b000_010001011100 : VALUE=19'b0000001_111010100111;
      15'b000_010001011101 : VALUE=19'b0000001_111010100100;
      15'b000_010001011110 : VALUE=19'b0000001_111010100000;
      15'b000_010001011111 : VALUE=19'b0000001_111010011101;
      15'b000_010001100000 : VALUE=19'b0000001_111010011001;
      15'b000_010001100001 : VALUE=19'b0000001_111010010110;
      15'b000_010001100010 : VALUE=19'b0000001_111010010010;
      15'b000_010001100011 : VALUE=19'b0000001_111010001111;
      15'b000_010001100100 : VALUE=19'b0000001_111010001011;
      15'b000_010001100101 : VALUE=19'b0000001_111010001000;
      15'b000_010001100110 : VALUE=19'b0000001_111010000100;
      15'b000_010001100111 : VALUE=19'b0000001_111010000001;
      15'b000_010001101000 : VALUE=19'b0000001_111001111101;
      15'b000_010001101001 : VALUE=19'b0000001_111001111010;
      15'b000_010001101010 : VALUE=19'b0000001_111001110110;
      15'b000_010001101011 : VALUE=19'b0000001_111001110011;
      15'b000_010001101100 : VALUE=19'b0000001_111001101111;
      15'b000_010001101101 : VALUE=19'b0000001_111001101100;
      15'b000_010001101110 : VALUE=19'b0000001_111001101001;
      15'b000_010001101111 : VALUE=19'b0000001_111001100101;
      15'b000_010001110000 : VALUE=19'b0000001_111001100010;
      15'b000_010001110001 : VALUE=19'b0000001_111001011110;
      15'b000_010001110010 : VALUE=19'b0000001_111001011011;
      15'b000_010001110011 : VALUE=19'b0000001_111001010111;
      15'b000_010001110100 : VALUE=19'b0000001_111001010100;
      15'b000_010001110101 : VALUE=19'b0000001_111001010001;
      15'b000_010001110110 : VALUE=19'b0000001_111001001101;
      15'b000_010001110111 : VALUE=19'b0000001_111001001010;
      15'b000_010001111000 : VALUE=19'b0000001_111001000110;
      15'b000_010001111001 : VALUE=19'b0000001_111001000011;
      15'b000_010001111010 : VALUE=19'b0000001_111001000000;
      15'b000_010001111011 : VALUE=19'b0000001_111000111100;
      15'b000_010001111100 : VALUE=19'b0000001_111000111001;
      15'b000_010001111101 : VALUE=19'b0000001_111000110110;
      15'b000_010001111110 : VALUE=19'b0000001_111000110010;
      15'b000_010001111111 : VALUE=19'b0000001_111000101111;
      15'b000_010010000000 : VALUE=19'b0000001_111000101011;
      15'b000_010010000001 : VALUE=19'b0000001_111000101000;
      15'b000_010010000010 : VALUE=19'b0000001_111000100101;
      15'b000_010010000011 : VALUE=19'b0000001_111000100001;
      15'b000_010010000100 : VALUE=19'b0000001_111000011110;
      15'b000_010010000101 : VALUE=19'b0000001_111000011011;
      15'b000_010010000110 : VALUE=19'b0000001_111000010111;
      15'b000_010010000111 : VALUE=19'b0000001_111000010100;
      15'b000_010010001000 : VALUE=19'b0000001_111000010001;
      15'b000_010010001001 : VALUE=19'b0000001_111000001101;
      15'b000_010010001010 : VALUE=19'b0000001_111000001010;
      15'b000_010010001011 : VALUE=19'b0000001_111000000111;
      15'b000_010010001100 : VALUE=19'b0000001_111000000100;
      15'b000_010010001101 : VALUE=19'b0000001_111000000000;
      15'b000_010010001110 : VALUE=19'b0000001_110111111101;
      15'b000_010010001111 : VALUE=19'b0000001_110111111010;
      15'b000_010010010000 : VALUE=19'b0000001_110111110110;
      15'b000_010010010001 : VALUE=19'b0000001_110111110011;
      15'b000_010010010010 : VALUE=19'b0000001_110111110000;
      15'b000_010010010011 : VALUE=19'b0000001_110111101101;
      15'b000_010010010100 : VALUE=19'b0000001_110111101001;
      15'b000_010010010101 : VALUE=19'b0000001_110111100110;
      15'b000_010010010110 : VALUE=19'b0000001_110111100011;
      15'b000_010010010111 : VALUE=19'b0000001_110111100000;
      15'b000_010010011000 : VALUE=19'b0000001_110111011100;
      15'b000_010010011001 : VALUE=19'b0000001_110111011001;
      15'b000_010010011010 : VALUE=19'b0000001_110111010110;
      15'b000_010010011011 : VALUE=19'b0000001_110111010011;
      15'b000_010010011100 : VALUE=19'b0000001_110111001111;
      15'b000_010010011101 : VALUE=19'b0000001_110111001100;
      15'b000_010010011110 : VALUE=19'b0000001_110111001001;
      15'b000_010010011111 : VALUE=19'b0000001_110111000110;
      15'b000_010010100000 : VALUE=19'b0000001_110111000010;
      15'b000_010010100001 : VALUE=19'b0000001_110110111111;
      15'b000_010010100010 : VALUE=19'b0000001_110110111100;
      15'b000_010010100011 : VALUE=19'b0000001_110110111001;
      15'b000_010010100100 : VALUE=19'b0000001_110110110110;
      15'b000_010010100101 : VALUE=19'b0000001_110110110010;
      15'b000_010010100110 : VALUE=19'b0000001_110110101111;
      15'b000_010010100111 : VALUE=19'b0000001_110110101100;
      15'b000_010010101000 : VALUE=19'b0000001_110110101001;
      15'b000_010010101001 : VALUE=19'b0000001_110110100110;
      15'b000_010010101010 : VALUE=19'b0000001_110110100010;
      15'b000_010010101011 : VALUE=19'b0000001_110110011111;
      15'b000_010010101100 : VALUE=19'b0000001_110110011100;
      15'b000_010010101101 : VALUE=19'b0000001_110110011001;
      15'b000_010010101110 : VALUE=19'b0000001_110110010110;
      15'b000_010010101111 : VALUE=19'b0000001_110110010011;
      15'b000_010010110000 : VALUE=19'b0000001_110110001111;
      15'b000_010010110001 : VALUE=19'b0000001_110110001100;
      15'b000_010010110010 : VALUE=19'b0000001_110110001001;
      15'b000_010010110011 : VALUE=19'b0000001_110110000110;
      15'b000_010010110100 : VALUE=19'b0000001_110110000011;
      15'b000_010010110101 : VALUE=19'b0000001_110110000000;
      15'b000_010010110110 : VALUE=19'b0000001_110101111101;
      15'b000_010010110111 : VALUE=19'b0000001_110101111001;
      15'b000_010010111000 : VALUE=19'b0000001_110101110110;
      15'b000_010010111001 : VALUE=19'b0000001_110101110011;
      15'b000_010010111010 : VALUE=19'b0000001_110101110000;
      15'b000_010010111011 : VALUE=19'b0000001_110101101101;
      15'b000_010010111100 : VALUE=19'b0000001_110101101010;
      15'b000_010010111101 : VALUE=19'b0000001_110101100111;
      15'b000_010010111110 : VALUE=19'b0000001_110101100100;
      15'b000_010010111111 : VALUE=19'b0000001_110101100001;
      15'b000_010011000000 : VALUE=19'b0000001_110101011101;
      15'b000_010011000001 : VALUE=19'b0000001_110101011010;
      15'b000_010011000010 : VALUE=19'b0000001_110101010111;
      15'b000_010011000011 : VALUE=19'b0000001_110101010100;
      15'b000_010011000100 : VALUE=19'b0000001_110101010001;
      15'b000_010011000101 : VALUE=19'b0000001_110101001110;
      15'b000_010011000110 : VALUE=19'b0000001_110101001011;
      15'b000_010011000111 : VALUE=19'b0000001_110101001000;
      15'b000_010011001000 : VALUE=19'b0000001_110101000101;
      15'b000_010011001001 : VALUE=19'b0000001_110101000010;
      15'b000_010011001010 : VALUE=19'b0000001_110100111111;
      15'b000_010011001011 : VALUE=19'b0000001_110100111100;
      15'b000_010011001100 : VALUE=19'b0000001_110100111001;
      15'b000_010011001101 : VALUE=19'b0000001_110100110110;
      15'b000_010011001110 : VALUE=19'b0000001_110100110011;
      15'b000_010011001111 : VALUE=19'b0000001_110100110000;
      15'b000_010011010000 : VALUE=19'b0000001_110100101101;
      15'b000_010011010001 : VALUE=19'b0000001_110100101001;
      15'b000_010011010010 : VALUE=19'b0000001_110100100110;
      15'b000_010011010011 : VALUE=19'b0000001_110100100011;
      15'b000_010011010100 : VALUE=19'b0000001_110100100000;
      15'b000_010011010101 : VALUE=19'b0000001_110100011101;
      15'b000_010011010110 : VALUE=19'b0000001_110100011010;
      15'b000_010011010111 : VALUE=19'b0000001_110100010111;
      15'b000_010011011000 : VALUE=19'b0000001_110100010100;
      15'b000_010011011001 : VALUE=19'b0000001_110100010001;
      15'b000_010011011010 : VALUE=19'b0000001_110100001110;
      15'b000_010011011011 : VALUE=19'b0000001_110100001011;
      15'b000_010011011100 : VALUE=19'b0000001_110100001000;
      15'b000_010011011101 : VALUE=19'b0000001_110100000101;
      15'b000_010011011110 : VALUE=19'b0000001_110100000010;
      15'b000_010011011111 : VALUE=19'b0000001_110011111111;
      15'b000_010011100000 : VALUE=19'b0000001_110011111100;
      15'b000_010011100001 : VALUE=19'b0000001_110011111010;
      15'b000_010011100010 : VALUE=19'b0000001_110011110111;
      15'b000_010011100011 : VALUE=19'b0000001_110011110100;
      15'b000_010011100100 : VALUE=19'b0000001_110011110001;
      15'b000_010011100101 : VALUE=19'b0000001_110011101110;
      15'b000_010011100110 : VALUE=19'b0000001_110011101011;
      15'b000_010011100111 : VALUE=19'b0000001_110011101000;
      15'b000_010011101000 : VALUE=19'b0000001_110011100101;
      15'b000_010011101001 : VALUE=19'b0000001_110011100010;
      15'b000_010011101010 : VALUE=19'b0000001_110011011111;
      15'b000_010011101011 : VALUE=19'b0000001_110011011100;
      15'b000_010011101100 : VALUE=19'b0000001_110011011001;
      15'b000_010011101101 : VALUE=19'b0000001_110011010110;
      15'b000_010011101110 : VALUE=19'b0000001_110011010011;
      15'b000_010011101111 : VALUE=19'b0000001_110011010000;
      15'b000_010011110000 : VALUE=19'b0000001_110011001101;
      15'b000_010011110001 : VALUE=19'b0000001_110011001010;
      15'b000_010011110010 : VALUE=19'b0000001_110011001000;
      15'b000_010011110011 : VALUE=19'b0000001_110011000101;
      15'b000_010011110100 : VALUE=19'b0000001_110011000010;
      15'b000_010011110101 : VALUE=19'b0000001_110010111111;
      15'b000_010011110110 : VALUE=19'b0000001_110010111100;
      15'b000_010011110111 : VALUE=19'b0000001_110010111001;
      15'b000_010011111000 : VALUE=19'b0000001_110010110110;
      15'b000_010011111001 : VALUE=19'b0000001_110010110011;
      15'b000_010011111010 : VALUE=19'b0000001_110010110000;
      15'b000_010011111011 : VALUE=19'b0000001_110010101110;
      15'b000_010011111100 : VALUE=19'b0000001_110010101011;
      15'b000_010011111101 : VALUE=19'b0000001_110010101000;
      15'b000_010011111110 : VALUE=19'b0000001_110010100101;
      15'b000_010011111111 : VALUE=19'b0000001_110010100010;
      15'b000_010100000000 : VALUE=19'b0000001_110010011111;
      15'b000_010100000001 : VALUE=19'b0000001_110010011100;
      15'b000_010100000010 : VALUE=19'b0000001_110010011001;
      15'b000_010100000011 : VALUE=19'b0000001_110010010111;
      15'b000_010100000100 : VALUE=19'b0000001_110010010100;
      15'b000_010100000101 : VALUE=19'b0000001_110010010001;
      15'b000_010100000110 : VALUE=19'b0000001_110010001110;
      15'b000_010100000111 : VALUE=19'b0000001_110010001011;
      15'b000_010100001000 : VALUE=19'b0000001_110010001000;
      15'b000_010100001001 : VALUE=19'b0000001_110010000110;
      15'b000_010100001010 : VALUE=19'b0000001_110010000011;
      15'b000_010100001011 : VALUE=19'b0000001_110010000000;
      15'b000_010100001100 : VALUE=19'b0000001_110001111101;
      15'b000_010100001101 : VALUE=19'b0000001_110001111010;
      15'b000_010100001110 : VALUE=19'b0000001_110001110111;
      15'b000_010100001111 : VALUE=19'b0000001_110001110101;
      15'b000_010100010000 : VALUE=19'b0000001_110001110010;
      15'b000_010100010001 : VALUE=19'b0000001_110001101111;
      15'b000_010100010010 : VALUE=19'b0000001_110001101100;
      15'b000_010100010011 : VALUE=19'b0000001_110001101001;
      15'b000_010100010100 : VALUE=19'b0000001_110001100111;
      15'b000_010100010101 : VALUE=19'b0000001_110001100100;
      15'b000_010100010110 : VALUE=19'b0000001_110001100001;
      15'b000_010100010111 : VALUE=19'b0000001_110001011110;
      15'b000_010100011000 : VALUE=19'b0000001_110001011011;
      15'b000_010100011001 : VALUE=19'b0000001_110001011001;
      15'b000_010100011010 : VALUE=19'b0000001_110001010110;
      15'b000_010100011011 : VALUE=19'b0000001_110001010011;
      15'b000_010100011100 : VALUE=19'b0000001_110001010000;
      15'b000_010100011101 : VALUE=19'b0000001_110001001110;
      15'b000_010100011110 : VALUE=19'b0000001_110001001011;
      15'b000_010100011111 : VALUE=19'b0000001_110001001000;
      15'b000_010100100000 : VALUE=19'b0000001_110001000101;
      15'b000_010100100001 : VALUE=19'b0000001_110001000010;
      15'b000_010100100010 : VALUE=19'b0000001_110001000000;
      15'b000_010100100011 : VALUE=19'b0000001_110000111101;
      15'b000_010100100100 : VALUE=19'b0000001_110000111010;
      15'b000_010100100101 : VALUE=19'b0000001_110000110111;
      15'b000_010100100110 : VALUE=19'b0000001_110000110101;
      15'b000_010100100111 : VALUE=19'b0000001_110000110010;
      15'b000_010100101000 : VALUE=19'b0000001_110000101111;
      15'b000_010100101001 : VALUE=19'b0000001_110000101101;
      15'b000_010100101010 : VALUE=19'b0000001_110000101010;
      15'b000_010100101011 : VALUE=19'b0000001_110000100111;
      15'b000_010100101100 : VALUE=19'b0000001_110000100100;
      15'b000_010100101101 : VALUE=19'b0000001_110000100010;
      15'b000_010100101110 : VALUE=19'b0000001_110000011111;
      15'b000_010100101111 : VALUE=19'b0000001_110000011100;
      15'b000_010100110000 : VALUE=19'b0000001_110000011010;
      15'b000_010100110001 : VALUE=19'b0000001_110000010111;
      15'b000_010100110010 : VALUE=19'b0000001_110000010100;
      15'b000_010100110011 : VALUE=19'b0000001_110000010001;
      15'b000_010100110100 : VALUE=19'b0000001_110000001111;
      15'b000_010100110101 : VALUE=19'b0000001_110000001100;
      15'b000_010100110110 : VALUE=19'b0000001_110000001001;
      15'b000_010100110111 : VALUE=19'b0000001_110000000111;
      15'b000_010100111000 : VALUE=19'b0000001_110000000100;
      15'b000_010100111001 : VALUE=19'b0000001_110000000001;
      15'b000_010100111010 : VALUE=19'b0000001_101111111111;
      15'b000_010100111011 : VALUE=19'b0000001_101111111100;
      15'b000_010100111100 : VALUE=19'b0000001_101111111001;
      15'b000_010100111101 : VALUE=19'b0000001_101111110111;
      15'b000_010100111110 : VALUE=19'b0000001_101111110100;
      15'b000_010100111111 : VALUE=19'b0000001_101111110001;
      15'b000_010101000000 : VALUE=19'b0000001_101111101111;
      15'b000_010101000001 : VALUE=19'b0000001_101111101100;
      15'b000_010101000010 : VALUE=19'b0000001_101111101001;
      15'b000_010101000011 : VALUE=19'b0000001_101111100111;
      15'b000_010101000100 : VALUE=19'b0000001_101111100100;
      15'b000_010101000101 : VALUE=19'b0000001_101111100001;
      15'b000_010101000110 : VALUE=19'b0000001_101111011111;
      15'b000_010101000111 : VALUE=19'b0000001_101111011100;
      15'b000_010101001000 : VALUE=19'b0000001_101111011001;
      15'b000_010101001001 : VALUE=19'b0000001_101111010111;
      15'b000_010101001010 : VALUE=19'b0000001_101111010100;
      15'b000_010101001011 : VALUE=19'b0000001_101111010001;
      15'b000_010101001100 : VALUE=19'b0000001_101111001111;
      15'b000_010101001101 : VALUE=19'b0000001_101111001100;
      15'b000_010101001110 : VALUE=19'b0000001_101111001010;
      15'b000_010101001111 : VALUE=19'b0000001_101111000111;
      15'b000_010101010000 : VALUE=19'b0000001_101111000100;
      15'b000_010101010001 : VALUE=19'b0000001_101111000010;
      15'b000_010101010010 : VALUE=19'b0000001_101110111111;
      15'b000_010101010011 : VALUE=19'b0000001_101110111101;
      15'b000_010101010100 : VALUE=19'b0000001_101110111010;
      15'b000_010101010101 : VALUE=19'b0000001_101110110111;
      15'b000_010101010110 : VALUE=19'b0000001_101110110101;
      15'b000_010101010111 : VALUE=19'b0000001_101110110010;
      15'b000_010101011000 : VALUE=19'b0000001_101110110000;
      15'b000_010101011001 : VALUE=19'b0000001_101110101101;
      15'b000_010101011010 : VALUE=19'b0000001_101110101010;
      15'b000_010101011011 : VALUE=19'b0000001_101110101000;
      15'b000_010101011100 : VALUE=19'b0000001_101110100101;
      15'b000_010101011101 : VALUE=19'b0000001_101110100011;
      15'b000_010101011110 : VALUE=19'b0000001_101110100000;
      15'b000_010101011111 : VALUE=19'b0000001_101110011101;
      15'b000_010101100000 : VALUE=19'b0000001_101110011011;
      15'b000_010101100001 : VALUE=19'b0000001_101110011000;
      15'b000_010101100010 : VALUE=19'b0000001_101110010110;
      15'b000_010101100011 : VALUE=19'b0000001_101110010011;
      15'b000_010101100100 : VALUE=19'b0000001_101110010001;
      15'b000_010101100101 : VALUE=19'b0000001_101110001110;
      15'b000_010101100110 : VALUE=19'b0000001_101110001100;
      15'b000_010101100111 : VALUE=19'b0000001_101110001001;
      15'b000_010101101000 : VALUE=19'b0000001_101110000110;
      15'b000_010101101001 : VALUE=19'b0000001_101110000100;
      15'b000_010101101010 : VALUE=19'b0000001_101110000001;
      15'b000_010101101011 : VALUE=19'b0000001_101101111111;
      15'b000_010101101100 : VALUE=19'b0000001_101101111100;
      15'b000_010101101101 : VALUE=19'b0000001_101101111010;
      15'b000_010101101110 : VALUE=19'b0000001_101101110111;
      15'b000_010101101111 : VALUE=19'b0000001_101101110101;
      15'b000_010101110000 : VALUE=19'b0000001_101101110010;
      15'b000_010101110001 : VALUE=19'b0000001_101101110000;
      15'b000_010101110010 : VALUE=19'b0000001_101101101101;
      15'b000_010101110011 : VALUE=19'b0000001_101101101011;
      15'b000_010101110100 : VALUE=19'b0000001_101101101000;
      15'b000_010101110101 : VALUE=19'b0000001_101101100110;
      15'b000_010101110110 : VALUE=19'b0000001_101101100011;
      15'b000_010101110111 : VALUE=19'b0000001_101101100001;
      15'b000_010101111000 : VALUE=19'b0000001_101101011110;
      15'b000_010101111001 : VALUE=19'b0000001_101101011100;
      15'b000_010101111010 : VALUE=19'b0000001_101101011001;
      15'b000_010101111011 : VALUE=19'b0000001_101101010111;
      15'b000_010101111100 : VALUE=19'b0000001_101101010100;
      15'b000_010101111101 : VALUE=19'b0000001_101101010010;
      15'b000_010101111110 : VALUE=19'b0000001_101101001111;
      15'b000_010101111111 : VALUE=19'b0000001_101101001101;
      15'b000_010110000000 : VALUE=19'b0000001_101101001010;
      15'b000_010110000001 : VALUE=19'b0000001_101101001000;
      15'b000_010110000010 : VALUE=19'b0000001_101101000101;
      15'b000_010110000011 : VALUE=19'b0000001_101101000011;
      15'b000_010110000100 : VALUE=19'b0000001_101101000000;
      15'b000_010110000101 : VALUE=19'b0000001_101100111110;
      15'b000_010110000110 : VALUE=19'b0000001_101100111011;
      15'b000_010110000111 : VALUE=19'b0000001_101100111001;
      15'b000_010110001000 : VALUE=19'b0000001_101100110110;
      15'b000_010110001001 : VALUE=19'b0000001_101100110100;
      15'b000_010110001010 : VALUE=19'b0000001_101100110001;
      15'b000_010110001011 : VALUE=19'b0000001_101100101111;
      15'b000_010110001100 : VALUE=19'b0000001_101100101101;
      15'b000_010110001101 : VALUE=19'b0000001_101100101010;
      15'b000_010110001110 : VALUE=19'b0000001_101100101000;
      15'b000_010110001111 : VALUE=19'b0000001_101100100101;
      15'b000_010110010000 : VALUE=19'b0000001_101100100011;
      15'b000_010110010001 : VALUE=19'b0000001_101100100000;
      15'b000_010110010010 : VALUE=19'b0000001_101100011110;
      15'b000_010110010011 : VALUE=19'b0000001_101100011011;
      15'b000_010110010100 : VALUE=19'b0000001_101100011001;
      15'b000_010110010101 : VALUE=19'b0000001_101100010111;
      15'b000_010110010110 : VALUE=19'b0000001_101100010100;
      15'b000_010110010111 : VALUE=19'b0000001_101100010010;
      15'b000_010110011000 : VALUE=19'b0000001_101100001111;
      15'b000_010110011001 : VALUE=19'b0000001_101100001101;
      15'b000_010110011010 : VALUE=19'b0000001_101100001011;
      15'b000_010110011011 : VALUE=19'b0000001_101100001000;
      15'b000_010110011100 : VALUE=19'b0000001_101100000110;
      15'b000_010110011101 : VALUE=19'b0000001_101100000011;
      15'b000_010110011110 : VALUE=19'b0000001_101100000001;
      15'b000_010110011111 : VALUE=19'b0000001_101011111111;
      15'b000_010110100000 : VALUE=19'b0000001_101011111100;
      15'b000_010110100001 : VALUE=19'b0000001_101011111010;
      15'b000_010110100010 : VALUE=19'b0000001_101011110111;
      15'b000_010110100011 : VALUE=19'b0000001_101011110101;
      15'b000_010110100100 : VALUE=19'b0000001_101011110011;
      15'b000_010110100101 : VALUE=19'b0000001_101011110000;
      15'b000_010110100110 : VALUE=19'b0000001_101011101110;
      15'b000_010110100111 : VALUE=19'b0000001_101011101011;
      15'b000_010110101000 : VALUE=19'b0000001_101011101001;
      15'b000_010110101001 : VALUE=19'b0000001_101011100111;
      15'b000_010110101010 : VALUE=19'b0000001_101011100100;
      15'b000_010110101011 : VALUE=19'b0000001_101011100010;
      15'b000_010110101100 : VALUE=19'b0000001_101011011111;
      15'b000_010110101101 : VALUE=19'b0000001_101011011101;
      15'b000_010110101110 : VALUE=19'b0000001_101011011011;
      15'b000_010110101111 : VALUE=19'b0000001_101011011000;
      15'b000_010110110000 : VALUE=19'b0000001_101011010110;
      15'b000_010110110001 : VALUE=19'b0000001_101011010100;
      15'b000_010110110010 : VALUE=19'b0000001_101011010001;
      15'b000_010110110011 : VALUE=19'b0000001_101011001111;
      15'b000_010110110100 : VALUE=19'b0000001_101011001101;
      15'b000_010110110101 : VALUE=19'b0000001_101011001010;
      15'b000_010110110110 : VALUE=19'b0000001_101011001000;
      15'b000_010110110111 : VALUE=19'b0000001_101011000110;
      15'b000_010110111000 : VALUE=19'b0000001_101011000011;
      15'b000_010110111001 : VALUE=19'b0000001_101011000001;
      15'b000_010110111010 : VALUE=19'b0000001_101010111111;
      15'b000_010110111011 : VALUE=19'b0000001_101010111100;
      15'b000_010110111100 : VALUE=19'b0000001_101010111010;
      15'b000_010110111101 : VALUE=19'b0000001_101010111000;
      15'b000_010110111110 : VALUE=19'b0000001_101010110101;
      15'b000_010110111111 : VALUE=19'b0000001_101010110011;
      15'b000_010111000000 : VALUE=19'b0000001_101010110001;
      15'b000_010111000001 : VALUE=19'b0000001_101010101110;
      15'b000_010111000010 : VALUE=19'b0000001_101010101100;
      15'b000_010111000011 : VALUE=19'b0000001_101010101010;
      15'b000_010111000100 : VALUE=19'b0000001_101010100111;
      15'b000_010111000101 : VALUE=19'b0000001_101010100101;
      15'b000_010111000110 : VALUE=19'b0000001_101010100011;
      15'b000_010111000111 : VALUE=19'b0000001_101010100000;
      15'b000_010111001000 : VALUE=19'b0000001_101010011110;
      15'b000_010111001001 : VALUE=19'b0000001_101010011100;
      15'b000_010111001010 : VALUE=19'b0000001_101010011010;
      15'b000_010111001011 : VALUE=19'b0000001_101010010111;
      15'b000_010111001100 : VALUE=19'b0000001_101010010101;
      15'b000_010111001101 : VALUE=19'b0000001_101010010011;
      15'b000_010111001110 : VALUE=19'b0000001_101010010000;
      15'b000_010111001111 : VALUE=19'b0000001_101010001110;
      15'b000_010111010000 : VALUE=19'b0000001_101010001100;
      15'b000_010111010001 : VALUE=19'b0000001_101010001001;
      15'b000_010111010010 : VALUE=19'b0000001_101010000111;
      15'b000_010111010011 : VALUE=19'b0000001_101010000101;
      15'b000_010111010100 : VALUE=19'b0000001_101010000011;
      15'b000_010111010101 : VALUE=19'b0000001_101010000000;
      15'b000_010111010110 : VALUE=19'b0000001_101001111110;
      15'b000_010111010111 : VALUE=19'b0000001_101001111100;
      15'b000_010111011000 : VALUE=19'b0000001_101001111010;
      15'b000_010111011001 : VALUE=19'b0000001_101001110111;
      15'b000_010111011010 : VALUE=19'b0000001_101001110101;
      15'b000_010111011011 : VALUE=19'b0000001_101001110011;
      15'b000_010111011100 : VALUE=19'b0000001_101001110001;
      15'b000_010111011101 : VALUE=19'b0000001_101001101110;
      15'b000_010111011110 : VALUE=19'b0000001_101001101100;
      15'b000_010111011111 : VALUE=19'b0000001_101001101010;
      15'b000_010111100000 : VALUE=19'b0000001_101001101000;
      15'b000_010111100001 : VALUE=19'b0000001_101001100101;
      15'b000_010111100010 : VALUE=19'b0000001_101001100011;
      15'b000_010111100011 : VALUE=19'b0000001_101001100001;
      15'b000_010111100100 : VALUE=19'b0000001_101001011111;
      15'b000_010111100101 : VALUE=19'b0000001_101001011100;
      15'b000_010111100110 : VALUE=19'b0000001_101001011010;
      15'b000_010111100111 : VALUE=19'b0000001_101001011000;
      15'b000_010111101000 : VALUE=19'b0000001_101001010110;
      15'b000_010111101001 : VALUE=19'b0000001_101001010011;
      15'b000_010111101010 : VALUE=19'b0000001_101001010001;
      15'b000_010111101011 : VALUE=19'b0000001_101001001111;
      15'b000_010111101100 : VALUE=19'b0000001_101001001101;
      15'b000_010111101101 : VALUE=19'b0000001_101001001010;
      15'b000_010111101110 : VALUE=19'b0000001_101001001000;
      15'b000_010111101111 : VALUE=19'b0000001_101001000110;
      15'b000_010111110000 : VALUE=19'b0000001_101001000100;
      15'b000_010111110001 : VALUE=19'b0000001_101001000010;
      15'b000_010111110010 : VALUE=19'b0000001_101000111111;
      15'b000_010111110011 : VALUE=19'b0000001_101000111101;
      15'b000_010111110100 : VALUE=19'b0000001_101000111011;
      15'b000_010111110101 : VALUE=19'b0000001_101000111001;
      15'b000_010111110110 : VALUE=19'b0000001_101000110111;
      15'b000_010111110111 : VALUE=19'b0000001_101000110100;
      15'b000_010111111000 : VALUE=19'b0000001_101000110010;
      15'b000_010111111001 : VALUE=19'b0000001_101000110000;
      15'b000_010111111010 : VALUE=19'b0000001_101000101110;
      15'b000_010111111011 : VALUE=19'b0000001_101000101100;
      15'b000_010111111100 : VALUE=19'b0000001_101000101001;
      15'b000_010111111101 : VALUE=19'b0000001_101000100111;
      15'b000_010111111110 : VALUE=19'b0000001_101000100101;
      15'b000_010111111111 : VALUE=19'b0000001_101000100011;
      15'b000_011000000000 : VALUE=19'b0000001_101000100001;
      15'b000_011000000001 : VALUE=19'b0000001_101000011111;
      15'b000_011000000010 : VALUE=19'b0000001_101000011100;
      15'b000_011000000011 : VALUE=19'b0000001_101000011010;
      15'b000_011000000100 : VALUE=19'b0000001_101000011000;
      15'b000_011000000101 : VALUE=19'b0000001_101000010110;
      15'b000_011000000110 : VALUE=19'b0000001_101000010100;
      15'b000_011000000111 : VALUE=19'b0000001_101000010010;
      15'b000_011000001000 : VALUE=19'b0000001_101000001111;
      15'b000_011000001001 : VALUE=19'b0000001_101000001101;
      15'b000_011000001010 : VALUE=19'b0000001_101000001011;
      15'b000_011000001011 : VALUE=19'b0000001_101000001001;
      15'b000_011000001100 : VALUE=19'b0000001_101000000111;
      15'b000_011000001101 : VALUE=19'b0000001_101000000101;
      15'b000_011000001110 : VALUE=19'b0000001_101000000010;
      15'b000_011000001111 : VALUE=19'b0000001_101000000000;
      15'b000_011000010000 : VALUE=19'b0000001_100111111110;
      15'b000_011000010001 : VALUE=19'b0000001_100111111100;
      15'b000_011000010010 : VALUE=19'b0000001_100111111010;
      15'b000_011000010011 : VALUE=19'b0000001_100111111000;
      15'b000_011000010100 : VALUE=19'b0000001_100111110110;
      15'b000_011000010101 : VALUE=19'b0000001_100111110011;
      15'b000_011000010110 : VALUE=19'b0000001_100111110001;
      15'b000_011000010111 : VALUE=19'b0000001_100111101111;
      15'b000_011000011000 : VALUE=19'b0000001_100111101101;
      15'b000_011000011001 : VALUE=19'b0000001_100111101011;
      15'b000_011000011010 : VALUE=19'b0000001_100111101001;
      15'b000_011000011011 : VALUE=19'b0000001_100111100111;
      15'b000_011000011100 : VALUE=19'b0000001_100111100101;
      15'b000_011000011101 : VALUE=19'b0000001_100111100010;
      15'b000_011000011110 : VALUE=19'b0000001_100111100000;
      15'b000_011000011111 : VALUE=19'b0000001_100111011110;
      15'b000_011000100000 : VALUE=19'b0000001_100111011100;
      15'b000_011000100001 : VALUE=19'b0000001_100111011010;
      15'b000_011000100010 : VALUE=19'b0000001_100111011000;
      15'b000_011000100011 : VALUE=19'b0000001_100111010110;
      15'b000_011000100100 : VALUE=19'b0000001_100111010100;
      15'b000_011000100101 : VALUE=19'b0000001_100111010010;
      15'b000_011000100110 : VALUE=19'b0000001_100111010000;
      15'b000_011000100111 : VALUE=19'b0000001_100111001101;
      15'b000_011000101000 : VALUE=19'b0000001_100111001011;
      15'b000_011000101001 : VALUE=19'b0000001_100111001001;
      15'b000_011000101010 : VALUE=19'b0000001_100111000111;
      15'b000_011000101011 : VALUE=19'b0000001_100111000101;
      15'b000_011000101100 : VALUE=19'b0000001_100111000011;
      15'b000_011000101101 : VALUE=19'b0000001_100111000001;
      15'b000_011000101110 : VALUE=19'b0000001_100110111111;
      15'b000_011000101111 : VALUE=19'b0000001_100110111101;
      15'b000_011000110000 : VALUE=19'b0000001_100110111011;
      15'b000_011000110001 : VALUE=19'b0000001_100110111001;
      15'b000_011000110010 : VALUE=19'b0000001_100110110110;
      15'b000_011000110011 : VALUE=19'b0000001_100110110100;
      15'b000_011000110100 : VALUE=19'b0000001_100110110010;
      15'b000_011000110101 : VALUE=19'b0000001_100110110000;
      15'b000_011000110110 : VALUE=19'b0000001_100110101110;
      15'b000_011000110111 : VALUE=19'b0000001_100110101100;
      15'b000_011000111000 : VALUE=19'b0000001_100110101010;
      15'b000_011000111001 : VALUE=19'b0000001_100110101000;
      15'b000_011000111010 : VALUE=19'b0000001_100110100110;
      15'b000_011000111011 : VALUE=19'b0000001_100110100100;
      15'b000_011000111100 : VALUE=19'b0000001_100110100010;
      15'b000_011000111101 : VALUE=19'b0000001_100110100000;
      15'b000_011000111110 : VALUE=19'b0000001_100110011110;
      15'b000_011000111111 : VALUE=19'b0000001_100110011100;
      15'b000_011001000000 : VALUE=19'b0000001_100110011010;
      15'b000_011001000001 : VALUE=19'b0000001_100110011000;
      15'b000_011001000010 : VALUE=19'b0000001_100110010110;
      15'b000_011001000011 : VALUE=19'b0000001_100110010011;
      15'b000_011001000100 : VALUE=19'b0000001_100110010001;
      15'b000_011001000101 : VALUE=19'b0000001_100110001111;
      15'b000_011001000110 : VALUE=19'b0000001_100110001101;
      15'b000_011001000111 : VALUE=19'b0000001_100110001011;
      15'b000_011001001000 : VALUE=19'b0000001_100110001001;
      15'b000_011001001001 : VALUE=19'b0000001_100110000111;
      15'b000_011001001010 : VALUE=19'b0000001_100110000101;
      15'b000_011001001011 : VALUE=19'b0000001_100110000011;
      15'b000_011001001100 : VALUE=19'b0000001_100110000001;
      15'b000_011001001101 : VALUE=19'b0000001_100101111111;
      15'b000_011001001110 : VALUE=19'b0000001_100101111101;
      15'b000_011001001111 : VALUE=19'b0000001_100101111011;
      15'b000_011001010000 : VALUE=19'b0000001_100101111001;
      15'b000_011001010001 : VALUE=19'b0000001_100101110111;
      15'b000_011001010010 : VALUE=19'b0000001_100101110101;
      15'b000_011001010011 : VALUE=19'b0000001_100101110011;
      15'b000_011001010100 : VALUE=19'b0000001_100101110001;
      15'b000_011001010101 : VALUE=19'b0000001_100101101111;
      15'b000_011001010110 : VALUE=19'b0000001_100101101101;
      15'b000_011001010111 : VALUE=19'b0000001_100101101011;
      15'b000_011001011000 : VALUE=19'b0000001_100101101001;
      15'b000_011001011001 : VALUE=19'b0000001_100101100111;
      15'b000_011001011010 : VALUE=19'b0000001_100101100101;
      15'b000_011001011011 : VALUE=19'b0000001_100101100011;
      15'b000_011001011100 : VALUE=19'b0000001_100101100001;
      15'b000_011001011101 : VALUE=19'b0000001_100101011111;
      15'b000_011001011110 : VALUE=19'b0000001_100101011101;
      15'b000_011001011111 : VALUE=19'b0000001_100101011011;
      15'b000_011001100000 : VALUE=19'b0000001_100101011001;
      15'b000_011001100001 : VALUE=19'b0000001_100101010111;
      15'b000_011001100010 : VALUE=19'b0000001_100101010101;
      15'b000_011001100011 : VALUE=19'b0000001_100101010011;
      15'b000_011001100100 : VALUE=19'b0000001_100101010001;
      15'b000_011001100101 : VALUE=19'b0000001_100101001111;
      15'b000_011001100110 : VALUE=19'b0000001_100101001101;
      15'b000_011001100111 : VALUE=19'b0000001_100101001011;
      15'b000_011001101000 : VALUE=19'b0000001_100101001001;
      15'b000_011001101001 : VALUE=19'b0000001_100101000111;
      15'b000_011001101010 : VALUE=19'b0000001_100101000101;
      15'b000_011001101011 : VALUE=19'b0000001_100101000011;
      15'b000_011001101100 : VALUE=19'b0000001_100101000001;
      15'b000_011001101101 : VALUE=19'b0000001_100100111111;
      15'b000_011001101110 : VALUE=19'b0000001_100100111101;
      15'b000_011001101111 : VALUE=19'b0000001_100100111011;
      15'b000_011001110000 : VALUE=19'b0000001_100100111001;
      15'b000_011001110001 : VALUE=19'b0000001_100100110111;
      15'b000_011001110010 : VALUE=19'b0000001_100100110110;
      15'b000_011001110011 : VALUE=19'b0000001_100100110100;
      15'b000_011001110100 : VALUE=19'b0000001_100100110010;
      15'b000_011001110101 : VALUE=19'b0000001_100100110000;
      15'b000_011001110110 : VALUE=19'b0000001_100100101110;
      15'b000_011001110111 : VALUE=19'b0000001_100100101100;
      15'b000_011001111000 : VALUE=19'b0000001_100100101010;
      15'b000_011001111001 : VALUE=19'b0000001_100100101000;
      15'b000_011001111010 : VALUE=19'b0000001_100100100110;
      15'b000_011001111011 : VALUE=19'b0000001_100100100100;
      15'b000_011001111100 : VALUE=19'b0000001_100100100010;
      15'b000_011001111101 : VALUE=19'b0000001_100100100000;
      15'b000_011001111110 : VALUE=19'b0000001_100100011110;
      15'b000_011001111111 : VALUE=19'b0000001_100100011100;
      15'b000_011010000000 : VALUE=19'b0000001_100100011010;
      15'b000_011010000001 : VALUE=19'b0000001_100100011000;
      15'b000_011010000010 : VALUE=19'b0000001_100100010110;
      15'b000_011010000011 : VALUE=19'b0000001_100100010101;
      15'b000_011010000100 : VALUE=19'b0000001_100100010011;
      15'b000_011010000101 : VALUE=19'b0000001_100100010001;
      15'b000_011010000110 : VALUE=19'b0000001_100100001111;
      15'b000_011010000111 : VALUE=19'b0000001_100100001101;
      15'b000_011010001000 : VALUE=19'b0000001_100100001011;
      15'b000_011010001001 : VALUE=19'b0000001_100100001001;
      15'b000_011010001010 : VALUE=19'b0000001_100100000111;
      15'b000_011010001011 : VALUE=19'b0000001_100100000101;
      15'b000_011010001100 : VALUE=19'b0000001_100100000011;
      15'b000_011010001101 : VALUE=19'b0000001_100100000001;
      15'b000_011010001110 : VALUE=19'b0000001_100011111111;
      15'b000_011010001111 : VALUE=19'b0000001_100011111110;
      15'b000_011010010000 : VALUE=19'b0000001_100011111100;
      15'b000_011010010001 : VALUE=19'b0000001_100011111010;
      15'b000_011010010010 : VALUE=19'b0000001_100011111000;
      15'b000_011010010011 : VALUE=19'b0000001_100011110110;
      15'b000_011010010100 : VALUE=19'b0000001_100011110100;
      15'b000_011010010101 : VALUE=19'b0000001_100011110010;
      15'b000_011010010110 : VALUE=19'b0000001_100011110000;
      15'b000_011010010111 : VALUE=19'b0000001_100011101110;
      15'b000_011010011000 : VALUE=19'b0000001_100011101100;
      15'b000_011010011001 : VALUE=19'b0000001_100011101011;
      15'b000_011010011010 : VALUE=19'b0000001_100011101001;
      15'b000_011010011011 : VALUE=19'b0000001_100011100111;
      15'b000_011010011100 : VALUE=19'b0000001_100011100101;
      15'b000_011010011101 : VALUE=19'b0000001_100011100011;
      15'b000_011010011110 : VALUE=19'b0000001_100011100001;
      15'b000_011010011111 : VALUE=19'b0000001_100011011111;
      15'b000_011010100000 : VALUE=19'b0000001_100011011101;
      15'b000_011010100001 : VALUE=19'b0000001_100011011100;
      15'b000_011010100010 : VALUE=19'b0000001_100011011010;
      15'b000_011010100011 : VALUE=19'b0000001_100011011000;
      15'b000_011010100100 : VALUE=19'b0000001_100011010110;
      15'b000_011010100101 : VALUE=19'b0000001_100011010100;
      15'b000_011010100110 : VALUE=19'b0000001_100011010010;
      15'b000_011010100111 : VALUE=19'b0000001_100011010000;
      15'b000_011010101000 : VALUE=19'b0000001_100011001110;
      15'b000_011010101001 : VALUE=19'b0000001_100011001101;
      15'b000_011010101010 : VALUE=19'b0000001_100011001011;
      15'b000_011010101011 : VALUE=19'b0000001_100011001001;
      15'b000_011010101100 : VALUE=19'b0000001_100011000111;
      15'b000_011010101101 : VALUE=19'b0000001_100011000101;
      15'b000_011010101110 : VALUE=19'b0000001_100011000011;
      15'b000_011010101111 : VALUE=19'b0000001_100011000001;
      15'b000_011010110000 : VALUE=19'b0000001_100011000000;
      15'b000_011010110001 : VALUE=19'b0000001_100010111110;
      15'b000_011010110010 : VALUE=19'b0000001_100010111100;
      15'b000_011010110011 : VALUE=19'b0000001_100010111010;
      15'b000_011010110100 : VALUE=19'b0000001_100010111000;
      15'b000_011010110101 : VALUE=19'b0000001_100010110110;
      15'b000_011010110110 : VALUE=19'b0000001_100010110101;
      15'b000_011010110111 : VALUE=19'b0000001_100010110011;
      15'b000_011010111000 : VALUE=19'b0000001_100010110001;
      15'b000_011010111001 : VALUE=19'b0000001_100010101111;
      15'b000_011010111010 : VALUE=19'b0000001_100010101101;
      15'b000_011010111011 : VALUE=19'b0000001_100010101011;
      15'b000_011010111100 : VALUE=19'b0000001_100010101010;
      15'b000_011010111101 : VALUE=19'b0000001_100010101000;
      15'b000_011010111110 : VALUE=19'b0000001_100010100110;
      15'b000_011010111111 : VALUE=19'b0000001_100010100100;
      15'b000_011011000000 : VALUE=19'b0000001_100010100010;
      15'b000_011011000001 : VALUE=19'b0000001_100010100000;
      15'b000_011011000010 : VALUE=19'b0000001_100010011111;
      15'b000_011011000011 : VALUE=19'b0000001_100010011101;
      15'b000_011011000100 : VALUE=19'b0000001_100010011011;
      15'b000_011011000101 : VALUE=19'b0000001_100010011001;
      15'b000_011011000110 : VALUE=19'b0000001_100010010111;
      15'b000_011011000111 : VALUE=19'b0000001_100010010101;
      15'b000_011011001000 : VALUE=19'b0000001_100010010100;
      15'b000_011011001001 : VALUE=19'b0000001_100010010010;
      15'b000_011011001010 : VALUE=19'b0000001_100010010000;
      15'b000_011011001011 : VALUE=19'b0000001_100010001110;
      15'b000_011011001100 : VALUE=19'b0000001_100010001100;
      15'b000_011011001101 : VALUE=19'b0000001_100010001011;
      15'b000_011011001110 : VALUE=19'b0000001_100010001001;
      15'b000_011011001111 : VALUE=19'b0000001_100010000111;
      15'b000_011011010000 : VALUE=19'b0000001_100010000101;
      15'b000_011011010001 : VALUE=19'b0000001_100010000011;
      15'b000_011011010010 : VALUE=19'b0000001_100010000010;
      15'b000_011011010011 : VALUE=19'b0000001_100010000000;
      15'b000_011011010100 : VALUE=19'b0000001_100001111110;
      15'b000_011011010101 : VALUE=19'b0000001_100001111100;
      15'b000_011011010110 : VALUE=19'b0000001_100001111010;
      15'b000_011011010111 : VALUE=19'b0000001_100001111001;
      15'b000_011011011000 : VALUE=19'b0000001_100001110111;
      15'b000_011011011001 : VALUE=19'b0000001_100001110101;
      15'b000_011011011010 : VALUE=19'b0000001_100001110011;
      15'b000_011011011011 : VALUE=19'b0000001_100001110010;
      15'b000_011011011100 : VALUE=19'b0000001_100001110000;
      15'b000_011011011101 : VALUE=19'b0000001_100001101110;
      15'b000_011011011110 : VALUE=19'b0000001_100001101100;
      15'b000_011011011111 : VALUE=19'b0000001_100001101010;
      15'b000_011011100000 : VALUE=19'b0000001_100001101001;
      15'b000_011011100001 : VALUE=19'b0000001_100001100111;
      15'b000_011011100010 : VALUE=19'b0000001_100001100101;
      15'b000_011011100011 : VALUE=19'b0000001_100001100011;
      15'b000_011011100100 : VALUE=19'b0000001_100001100010;
      15'b000_011011100101 : VALUE=19'b0000001_100001100000;
      15'b000_011011100110 : VALUE=19'b0000001_100001011110;
      15'b000_011011100111 : VALUE=19'b0000001_100001011100;
      15'b000_011011101000 : VALUE=19'b0000001_100001011010;
      15'b000_011011101001 : VALUE=19'b0000001_100001011001;
      15'b000_011011101010 : VALUE=19'b0000001_100001010111;
      15'b000_011011101011 : VALUE=19'b0000001_100001010101;
      15'b000_011011101100 : VALUE=19'b0000001_100001010011;
      15'b000_011011101101 : VALUE=19'b0000001_100001010010;
      15'b000_011011101110 : VALUE=19'b0000001_100001010000;
      15'b000_011011101111 : VALUE=19'b0000001_100001001110;
      15'b000_011011110000 : VALUE=19'b0000001_100001001100;
      15'b000_011011110001 : VALUE=19'b0000001_100001001011;
      15'b000_011011110010 : VALUE=19'b0000001_100001001001;
      15'b000_011011110011 : VALUE=19'b0000001_100001000111;
      15'b000_011011110100 : VALUE=19'b0000001_100001000101;
      15'b000_011011110101 : VALUE=19'b0000001_100001000100;
      15'b000_011011110110 : VALUE=19'b0000001_100001000010;
      15'b000_011011110111 : VALUE=19'b0000001_100001000000;
      15'b000_011011111000 : VALUE=19'b0000001_100000111110;
      15'b000_011011111001 : VALUE=19'b0000001_100000111101;
      15'b000_011011111010 : VALUE=19'b0000001_100000111011;
      15'b000_011011111011 : VALUE=19'b0000001_100000111001;
      15'b000_011011111100 : VALUE=19'b0000001_100000110111;
      15'b000_011011111101 : VALUE=19'b0000001_100000110110;
      15'b000_011011111110 : VALUE=19'b0000001_100000110100;
      15'b000_011011111111 : VALUE=19'b0000001_100000110010;
      15'b000_011100000000 : VALUE=19'b0000001_100000110001;
      15'b000_011100000001 : VALUE=19'b0000001_100000101111;
      15'b000_011100000010 : VALUE=19'b0000001_100000101101;
      15'b000_011100000011 : VALUE=19'b0000001_100000101011;
      15'b000_011100000100 : VALUE=19'b0000001_100000101010;
      15'b000_011100000101 : VALUE=19'b0000001_100000101000;
      15'b000_011100000110 : VALUE=19'b0000001_100000100110;
      15'b000_011100000111 : VALUE=19'b0000001_100000100101;
      15'b000_011100001000 : VALUE=19'b0000001_100000100011;
      15'b000_011100001001 : VALUE=19'b0000001_100000100001;
      15'b000_011100001010 : VALUE=19'b0000001_100000011111;
      15'b000_011100001011 : VALUE=19'b0000001_100000011110;
      15'b000_011100001100 : VALUE=19'b0000001_100000011100;
      15'b000_011100001101 : VALUE=19'b0000001_100000011010;
      15'b000_011100001110 : VALUE=19'b0000001_100000011001;
      15'b000_011100001111 : VALUE=19'b0000001_100000010111;
      15'b000_011100010000 : VALUE=19'b0000001_100000010101;
      15'b000_011100010001 : VALUE=19'b0000001_100000010011;
      15'b000_011100010010 : VALUE=19'b0000001_100000010010;
      15'b000_011100010011 : VALUE=19'b0000001_100000010000;
      15'b000_011100010100 : VALUE=19'b0000001_100000001110;
      15'b000_011100010101 : VALUE=19'b0000001_100000001101;
      15'b000_011100010110 : VALUE=19'b0000001_100000001011;
      15'b000_011100010111 : VALUE=19'b0000001_100000001001;
      15'b000_011100011000 : VALUE=19'b0000001_100000001000;
      15'b000_011100011001 : VALUE=19'b0000001_100000000110;
      15'b000_011100011010 : VALUE=19'b0000001_100000000100;
      15'b000_011100011011 : VALUE=19'b0000001_100000000010;
      15'b000_011100011100 : VALUE=19'b0000001_100000000001;
      15'b000_011100011101 : VALUE=19'b0000001_011111111111;
      15'b000_011100011110 : VALUE=19'b0000001_011111111101;
      15'b000_011100011111 : VALUE=19'b0000001_011111111100;
      15'b000_011100100000 : VALUE=19'b0000001_011111111010;
      15'b000_011100100001 : VALUE=19'b0000001_011111111000;
      15'b000_011100100010 : VALUE=19'b0000001_011111110111;
      15'b000_011100100011 : VALUE=19'b0000001_011111110101;
      15'b000_011100100100 : VALUE=19'b0000001_011111110011;
      15'b000_011100100101 : VALUE=19'b0000001_011111110010;
      15'b000_011100100110 : VALUE=19'b0000001_011111110000;
      15'b000_011100100111 : VALUE=19'b0000001_011111101110;
      15'b000_011100101000 : VALUE=19'b0000001_011111101101;
      15'b000_011100101001 : VALUE=19'b0000001_011111101011;
      15'b000_011100101010 : VALUE=19'b0000001_011111101001;
      15'b000_011100101011 : VALUE=19'b0000001_011111101000;
      15'b000_011100101100 : VALUE=19'b0000001_011111100110;
      15'b000_011100101101 : VALUE=19'b0000001_011111100100;
      15'b000_011100101110 : VALUE=19'b0000001_011111100011;
      15'b000_011100101111 : VALUE=19'b0000001_011111100001;
      15'b000_011100110000 : VALUE=19'b0000001_011111011111;
      15'b000_011100110001 : VALUE=19'b0000001_011111011110;
      15'b000_011100110010 : VALUE=19'b0000001_011111011100;
      15'b000_011100110011 : VALUE=19'b0000001_011111011010;
      15'b000_011100110100 : VALUE=19'b0000001_011111011001;
      15'b000_011100110101 : VALUE=19'b0000001_011111010111;
      15'b000_011100110110 : VALUE=19'b0000001_011111010101;
      15'b000_011100110111 : VALUE=19'b0000001_011111010100;
      15'b000_011100111000 : VALUE=19'b0000001_011111010010;
      15'b000_011100111001 : VALUE=19'b0000001_011111010000;
      15'b000_011100111010 : VALUE=19'b0000001_011111001111;
      15'b000_011100111011 : VALUE=19'b0000001_011111001101;
      15'b000_011100111100 : VALUE=19'b0000001_011111001011;
      15'b000_011100111101 : VALUE=19'b0000001_011111001010;
      15'b000_011100111110 : VALUE=19'b0000001_011111001000;
      15'b000_011100111111 : VALUE=19'b0000001_011111000111;
      15'b000_011101000000 : VALUE=19'b0000001_011111000101;
      15'b000_011101000001 : VALUE=19'b0000001_011111000011;
      15'b000_011101000010 : VALUE=19'b0000001_011111000010;
      15'b000_011101000011 : VALUE=19'b0000001_011111000000;
      15'b000_011101000100 : VALUE=19'b0000001_011110111110;
      15'b000_011101000101 : VALUE=19'b0000001_011110111101;
      15'b000_011101000110 : VALUE=19'b0000001_011110111011;
      15'b000_011101000111 : VALUE=19'b0000001_011110111001;
      15'b000_011101001000 : VALUE=19'b0000001_011110111000;
      15'b000_011101001001 : VALUE=19'b0000001_011110110110;
      15'b000_011101001010 : VALUE=19'b0000001_011110110101;
      15'b000_011101001011 : VALUE=19'b0000001_011110110011;
      15'b000_011101001100 : VALUE=19'b0000001_011110110001;
      15'b000_011101001101 : VALUE=19'b0000001_011110110000;
      15'b000_011101001110 : VALUE=19'b0000001_011110101110;
      15'b000_011101001111 : VALUE=19'b0000001_011110101100;
      15'b000_011101010000 : VALUE=19'b0000001_011110101011;
      15'b000_011101010001 : VALUE=19'b0000001_011110101001;
      15'b000_011101010010 : VALUE=19'b0000001_011110101000;
      15'b000_011101010011 : VALUE=19'b0000001_011110100110;
      15'b000_011101010100 : VALUE=19'b0000001_011110100100;
      15'b000_011101010101 : VALUE=19'b0000001_011110100011;
      15'b000_011101010110 : VALUE=19'b0000001_011110100001;
      15'b000_011101010111 : VALUE=19'b0000001_011110100000;
      15'b000_011101011000 : VALUE=19'b0000001_011110011110;
      15'b000_011101011001 : VALUE=19'b0000001_011110011100;
      15'b000_011101011010 : VALUE=19'b0000001_011110011011;
      15'b000_011101011011 : VALUE=19'b0000001_011110011001;
      15'b000_011101011100 : VALUE=19'b0000001_011110010111;
      15'b000_011101011101 : VALUE=19'b0000001_011110010110;
      15'b000_011101011110 : VALUE=19'b0000001_011110010100;
      15'b000_011101011111 : VALUE=19'b0000001_011110010011;
      15'b000_011101100000 : VALUE=19'b0000001_011110010001;
      15'b000_011101100001 : VALUE=19'b0000001_011110001111;
      15'b000_011101100010 : VALUE=19'b0000001_011110001110;
      15'b000_011101100011 : VALUE=19'b0000001_011110001100;
      15'b000_011101100100 : VALUE=19'b0000001_011110001011;
      15'b000_011101100101 : VALUE=19'b0000001_011110001001;
      15'b000_011101100110 : VALUE=19'b0000001_011110001000;
      15'b000_011101100111 : VALUE=19'b0000001_011110000110;
      15'b000_011101101000 : VALUE=19'b0000001_011110000100;
      15'b000_011101101001 : VALUE=19'b0000001_011110000011;
      15'b000_011101101010 : VALUE=19'b0000001_011110000001;
      15'b000_011101101011 : VALUE=19'b0000001_011110000000;
      15'b000_011101101100 : VALUE=19'b0000001_011101111110;
      15'b000_011101101101 : VALUE=19'b0000001_011101111100;
      15'b000_011101101110 : VALUE=19'b0000001_011101111011;
      15'b000_011101101111 : VALUE=19'b0000001_011101111001;
      15'b000_011101110000 : VALUE=19'b0000001_011101111000;
      15'b000_011101110001 : VALUE=19'b0000001_011101110110;
      15'b000_011101110010 : VALUE=19'b0000001_011101110101;
      15'b000_011101110011 : VALUE=19'b0000001_011101110011;
      15'b000_011101110100 : VALUE=19'b0000001_011101110001;
      15'b000_011101110101 : VALUE=19'b0000001_011101110000;
      15'b000_011101110110 : VALUE=19'b0000001_011101101110;
      15'b000_011101110111 : VALUE=19'b0000001_011101101101;
      15'b000_011101111000 : VALUE=19'b0000001_011101101011;
      15'b000_011101111001 : VALUE=19'b0000001_011101101010;
      15'b000_011101111010 : VALUE=19'b0000001_011101101000;
      15'b000_011101111011 : VALUE=19'b0000001_011101100110;
      15'b000_011101111100 : VALUE=19'b0000001_011101100101;
      15'b000_011101111101 : VALUE=19'b0000001_011101100011;
      15'b000_011101111110 : VALUE=19'b0000001_011101100010;
      15'b000_011101111111 : VALUE=19'b0000001_011101100000;
      15'b000_011110000000 : VALUE=19'b0000001_011101011111;
      15'b000_011110000001 : VALUE=19'b0000001_011101011101;
      15'b000_011110000010 : VALUE=19'b0000001_011101011011;
      15'b000_011110000011 : VALUE=19'b0000001_011101011010;
      15'b000_011110000100 : VALUE=19'b0000001_011101011000;
      15'b000_011110000101 : VALUE=19'b0000001_011101010111;
      15'b000_011110000110 : VALUE=19'b0000001_011101010101;
      15'b000_011110000111 : VALUE=19'b0000001_011101010100;
      15'b000_011110001000 : VALUE=19'b0000001_011101010010;
      15'b000_011110001001 : VALUE=19'b0000001_011101010001;
      15'b000_011110001010 : VALUE=19'b0000001_011101001111;
      15'b000_011110001011 : VALUE=19'b0000001_011101001110;
      15'b000_011110001100 : VALUE=19'b0000001_011101001100;
      15'b000_011110001101 : VALUE=19'b0000001_011101001010;
      15'b000_011110001110 : VALUE=19'b0000001_011101001001;
      15'b000_011110001111 : VALUE=19'b0000001_011101000111;
      15'b000_011110010000 : VALUE=19'b0000001_011101000110;
      15'b000_011110010001 : VALUE=19'b0000001_011101000100;
      15'b000_011110010010 : VALUE=19'b0000001_011101000011;
      15'b000_011110010011 : VALUE=19'b0000001_011101000001;
      15'b000_011110010100 : VALUE=19'b0000001_011101000000;
      15'b000_011110010101 : VALUE=19'b0000001_011100111110;
      15'b000_011110010110 : VALUE=19'b0000001_011100111101;
      15'b000_011110010111 : VALUE=19'b0000001_011100111011;
      15'b000_011110011000 : VALUE=19'b0000001_011100111010;
      15'b000_011110011001 : VALUE=19'b0000001_011100111000;
      15'b000_011110011010 : VALUE=19'b0000001_011100110110;
      15'b000_011110011011 : VALUE=19'b0000001_011100110101;
      15'b000_011110011100 : VALUE=19'b0000001_011100110011;
      15'b000_011110011101 : VALUE=19'b0000001_011100110010;
      15'b000_011110011110 : VALUE=19'b0000001_011100110000;
      15'b000_011110011111 : VALUE=19'b0000001_011100101111;
      15'b000_011110100000 : VALUE=19'b0000001_011100101101;
      15'b000_011110100001 : VALUE=19'b0000001_011100101100;
      15'b000_011110100010 : VALUE=19'b0000001_011100101010;
      15'b000_011110100011 : VALUE=19'b0000001_011100101001;
      15'b000_011110100100 : VALUE=19'b0000001_011100100111;
      15'b000_011110100101 : VALUE=19'b0000001_011100100110;
      15'b000_011110100110 : VALUE=19'b0000001_011100100100;
      15'b000_011110100111 : VALUE=19'b0000001_011100100011;
      15'b000_011110101000 : VALUE=19'b0000001_011100100001;
      15'b000_011110101001 : VALUE=19'b0000001_011100100000;
      15'b000_011110101010 : VALUE=19'b0000001_011100011110;
      15'b000_011110101011 : VALUE=19'b0000001_011100011101;
      15'b000_011110101100 : VALUE=19'b0000001_011100011011;
      15'b000_011110101101 : VALUE=19'b0000001_011100011010;
      15'b000_011110101110 : VALUE=19'b0000001_011100011000;
      15'b000_011110101111 : VALUE=19'b0000001_011100010111;
      15'b000_011110110000 : VALUE=19'b0000001_011100010101;
      15'b000_011110110001 : VALUE=19'b0000001_011100010100;
      15'b000_011110110010 : VALUE=19'b0000001_011100010010;
      15'b000_011110110011 : VALUE=19'b0000001_011100010001;
      15'b000_011110110100 : VALUE=19'b0000001_011100001111;
      15'b000_011110110101 : VALUE=19'b0000001_011100001110;
      15'b000_011110110110 : VALUE=19'b0000001_011100001100;
      15'b000_011110110111 : VALUE=19'b0000001_011100001011;
      15'b000_011110111000 : VALUE=19'b0000001_011100001001;
      15'b000_011110111001 : VALUE=19'b0000001_011100001000;
      15'b000_011110111010 : VALUE=19'b0000001_011100000110;
      15'b000_011110111011 : VALUE=19'b0000001_011100000101;
      15'b000_011110111100 : VALUE=19'b0000001_011100000011;
      15'b000_011110111101 : VALUE=19'b0000001_011100000010;
      15'b000_011110111110 : VALUE=19'b0000001_011100000000;
      15'b000_011110111111 : VALUE=19'b0000001_011011111111;
      15'b000_011111000000 : VALUE=19'b0000001_011011111101;
      15'b000_011111000001 : VALUE=19'b0000001_011011111100;
      15'b000_011111000010 : VALUE=19'b0000001_011011111010;
      15'b000_011111000011 : VALUE=19'b0000001_011011111001;
      15'b000_011111000100 : VALUE=19'b0000001_011011110111;
      15'b000_011111000101 : VALUE=19'b0000001_011011110110;
      15'b000_011111000110 : VALUE=19'b0000001_011011110100;
      15'b000_011111000111 : VALUE=19'b0000001_011011110011;
      15'b000_011111001000 : VALUE=19'b0000001_011011110001;
      15'b000_011111001001 : VALUE=19'b0000001_011011110000;
      15'b000_011111001010 : VALUE=19'b0000001_011011101111;
      15'b000_011111001011 : VALUE=19'b0000001_011011101101;
      15'b000_011111001100 : VALUE=19'b0000001_011011101100;
      15'b000_011111001101 : VALUE=19'b0000001_011011101010;
      15'b000_011111001110 : VALUE=19'b0000001_011011101001;
      15'b000_011111001111 : VALUE=19'b0000001_011011100111;
      15'b000_011111010000 : VALUE=19'b0000001_011011100110;
      15'b000_011111010001 : VALUE=19'b0000001_011011100100;
      15'b000_011111010010 : VALUE=19'b0000001_011011100011;
      15'b000_011111010011 : VALUE=19'b0000001_011011100001;
      15'b000_011111010100 : VALUE=19'b0000001_011011100000;
      15'b000_011111010101 : VALUE=19'b0000001_011011011110;
      15'b000_011111010110 : VALUE=19'b0000001_011011011101;
      15'b000_011111010111 : VALUE=19'b0000001_011011011011;
      15'b000_011111011000 : VALUE=19'b0000001_011011011010;
      15'b000_011111011001 : VALUE=19'b0000001_011011011001;
      15'b000_011111011010 : VALUE=19'b0000001_011011010111;
      15'b000_011111011011 : VALUE=19'b0000001_011011010110;
      15'b000_011111011100 : VALUE=19'b0000001_011011010100;
      15'b000_011111011101 : VALUE=19'b0000001_011011010011;
      15'b000_011111011110 : VALUE=19'b0000001_011011010001;
      15'b000_011111011111 : VALUE=19'b0000001_011011010000;
      15'b000_011111100000 : VALUE=19'b0000001_011011001110;
      15'b000_011111100001 : VALUE=19'b0000001_011011001101;
      15'b000_011111100010 : VALUE=19'b0000001_011011001100;
      15'b000_011111100011 : VALUE=19'b0000001_011011001010;
      15'b000_011111100100 : VALUE=19'b0000001_011011001001;
      15'b000_011111100101 : VALUE=19'b0000001_011011000111;
      15'b000_011111100110 : VALUE=19'b0000001_011011000110;
      15'b000_011111100111 : VALUE=19'b0000001_011011000100;
      15'b000_011111101000 : VALUE=19'b0000001_011011000011;
      15'b000_011111101001 : VALUE=19'b0000001_011011000001;
      15'b000_011111101010 : VALUE=19'b0000001_011011000000;
      15'b000_011111101011 : VALUE=19'b0000001_011010111111;
      15'b000_011111101100 : VALUE=19'b0000001_011010111101;
      15'b000_011111101101 : VALUE=19'b0000001_011010111100;
      15'b000_011111101110 : VALUE=19'b0000001_011010111010;
      15'b000_011111101111 : VALUE=19'b0000001_011010111001;
      15'b000_011111110000 : VALUE=19'b0000001_011010110111;
      15'b000_011111110001 : VALUE=19'b0000001_011010110110;
      15'b000_011111110010 : VALUE=19'b0000001_011010110101;
      15'b000_011111110011 : VALUE=19'b0000001_011010110011;
      15'b000_011111110100 : VALUE=19'b0000001_011010110010;
      15'b000_011111110101 : VALUE=19'b0000001_011010110000;
      15'b000_011111110110 : VALUE=19'b0000001_011010101111;
      15'b000_011111110111 : VALUE=19'b0000001_011010101101;
      15'b000_011111111000 : VALUE=19'b0000001_011010101100;
      15'b000_011111111001 : VALUE=19'b0000001_011010101011;
      15'b000_011111111010 : VALUE=19'b0000001_011010101001;
      15'b000_011111111011 : VALUE=19'b0000001_011010101000;
      15'b000_011111111100 : VALUE=19'b0000001_011010100110;
      15'b000_011111111101 : VALUE=19'b0000001_011010100101;
      15'b000_011111111110 : VALUE=19'b0000001_011010100011;
      15'b000_011111111111 : VALUE=19'b0000001_011010100010;
      15'b000_100000000000 : VALUE=19'b0000001_011010100001;
      15'b000_100000000001 : VALUE=19'b0000001_011010011111;
      15'b000_100000000010 : VALUE=19'b0000001_011010011110;
      15'b000_100000000011 : VALUE=19'b0000001_011010011100;
      15'b000_100000000100 : VALUE=19'b0000001_011010011011;
      15'b000_100000000101 : VALUE=19'b0000001_011010011010;
      15'b000_100000000110 : VALUE=19'b0000001_011010011000;
      15'b000_100000000111 : VALUE=19'b0000001_011010010111;
      15'b000_100000001000 : VALUE=19'b0000001_011010010101;
      15'b000_100000001001 : VALUE=19'b0000001_011010010100;
      15'b000_100000001010 : VALUE=19'b0000001_011010010011;
      15'b000_100000001011 : VALUE=19'b0000001_011010010001;
      15'b000_100000001100 : VALUE=19'b0000001_011010010000;
      15'b000_100000001101 : VALUE=19'b0000001_011010001110;
      15'b000_100000001110 : VALUE=19'b0000001_011010001101;
      15'b000_100000001111 : VALUE=19'b0000001_011010001100;
      15'b000_100000010000 : VALUE=19'b0000001_011010001010;
      15'b000_100000010001 : VALUE=19'b0000001_011010001001;
      15'b000_100000010010 : VALUE=19'b0000001_011010000111;
      15'b000_100000010011 : VALUE=19'b0000001_011010000110;
      15'b000_100000010100 : VALUE=19'b0000001_011010000101;
      15'b000_100000010101 : VALUE=19'b0000001_011010000011;
      15'b000_100000010110 : VALUE=19'b0000001_011010000010;
      15'b000_100000010111 : VALUE=19'b0000001_011010000000;
      15'b000_100000011000 : VALUE=19'b0000001_011001111111;
      15'b000_100000011001 : VALUE=19'b0000001_011001111110;
      15'b000_100000011010 : VALUE=19'b0000001_011001111100;
      15'b000_100000011011 : VALUE=19'b0000001_011001111011;
      15'b000_100000011100 : VALUE=19'b0000001_011001111001;
      15'b000_100000011101 : VALUE=19'b0000001_011001111000;
      15'b000_100000011110 : VALUE=19'b0000001_011001110111;
      15'b000_100000011111 : VALUE=19'b0000001_011001110101;
      15'b000_100000100000 : VALUE=19'b0000001_011001110100;
      15'b000_100000100001 : VALUE=19'b0000001_011001110011;
      15'b000_100000100010 : VALUE=19'b0000001_011001110001;
      15'b000_100000100011 : VALUE=19'b0000001_011001110000;
      15'b000_100000100100 : VALUE=19'b0000001_011001101110;
      15'b000_100000100101 : VALUE=19'b0000001_011001101101;
      15'b000_100000100110 : VALUE=19'b0000001_011001101100;
      15'b000_100000100111 : VALUE=19'b0000001_011001101010;
      15'b000_100000101000 : VALUE=19'b0000001_011001101001;
      15'b000_100000101001 : VALUE=19'b0000001_011001100111;
      15'b000_100000101010 : VALUE=19'b0000001_011001100110;
      15'b000_100000101011 : VALUE=19'b0000001_011001100101;
      15'b000_100000101100 : VALUE=19'b0000001_011001100011;
      15'b000_100000101101 : VALUE=19'b0000001_011001100010;
      15'b000_100000101110 : VALUE=19'b0000001_011001100001;
      15'b000_100000101111 : VALUE=19'b0000001_011001011111;
      15'b000_100000110000 : VALUE=19'b0000001_011001011110;
      15'b000_100000110001 : VALUE=19'b0000001_011001011101;
      15'b000_100000110010 : VALUE=19'b0000001_011001011011;
      15'b000_100000110011 : VALUE=19'b0000001_011001011010;
      15'b000_100000110100 : VALUE=19'b0000001_011001011000;
      15'b000_100000110101 : VALUE=19'b0000001_011001010111;
      15'b000_100000110110 : VALUE=19'b0000001_011001010110;
      15'b000_100000110111 : VALUE=19'b0000001_011001010100;
      15'b000_100000111000 : VALUE=19'b0000001_011001010011;
      15'b000_100000111001 : VALUE=19'b0000001_011001010010;
      15'b000_100000111010 : VALUE=19'b0000001_011001010000;
      15'b000_100000111011 : VALUE=19'b0000001_011001001111;
      15'b000_100000111100 : VALUE=19'b0000001_011001001110;
      15'b000_100000111101 : VALUE=19'b0000001_011001001100;
      15'b000_100000111110 : VALUE=19'b0000001_011001001011;
      15'b000_100000111111 : VALUE=19'b0000001_011001001010;
      15'b000_100001000000 : VALUE=19'b0000001_011001001000;
      15'b000_100001000001 : VALUE=19'b0000001_011001000111;
      15'b000_100001000010 : VALUE=19'b0000001_011001000101;
      15'b000_100001000011 : VALUE=19'b0000001_011001000100;
      15'b000_100001000100 : VALUE=19'b0000001_011001000011;
      15'b000_100001000101 : VALUE=19'b0000001_011001000001;
      15'b000_100001000110 : VALUE=19'b0000001_011001000000;
      15'b000_100001000111 : VALUE=19'b0000001_011000111111;
      15'b000_100001001000 : VALUE=19'b0000001_011000111101;
      15'b000_100001001001 : VALUE=19'b0000001_011000111100;
      15'b000_100001001010 : VALUE=19'b0000001_011000111011;
      15'b000_100001001011 : VALUE=19'b0000001_011000111001;
      15'b000_100001001100 : VALUE=19'b0000001_011000111000;
      15'b000_100001001101 : VALUE=19'b0000001_011000110111;
      15'b000_100001001110 : VALUE=19'b0000001_011000110101;
      15'b000_100001001111 : VALUE=19'b0000001_011000110100;
      15'b000_100001010000 : VALUE=19'b0000001_011000110011;
      15'b000_100001010001 : VALUE=19'b0000001_011000110001;
      15'b000_100001010010 : VALUE=19'b0000001_011000110000;
      15'b000_100001010011 : VALUE=19'b0000001_011000101111;
      15'b000_100001010100 : VALUE=19'b0000001_011000101101;
      15'b000_100001010101 : VALUE=19'b0000001_011000101100;
      15'b000_100001010110 : VALUE=19'b0000001_011000101011;
      15'b000_100001010111 : VALUE=19'b0000001_011000101001;
      15'b000_100001011000 : VALUE=19'b0000001_011000101000;
      15'b000_100001011001 : VALUE=19'b0000001_011000100111;
      15'b000_100001011010 : VALUE=19'b0000001_011000100101;
      15'b000_100001011011 : VALUE=19'b0000001_011000100100;
      15'b000_100001011100 : VALUE=19'b0000001_011000100011;
      15'b000_100001011101 : VALUE=19'b0000001_011000100001;
      15'b000_100001011110 : VALUE=19'b0000001_011000100000;
      15'b000_100001011111 : VALUE=19'b0000001_011000011111;
      15'b000_100001100000 : VALUE=19'b0000001_011000011101;
      15'b000_100001100001 : VALUE=19'b0000001_011000011100;
      15'b000_100001100010 : VALUE=19'b0000001_011000011011;
      15'b000_100001100011 : VALUE=19'b0000001_011000011001;
      15'b000_100001100100 : VALUE=19'b0000001_011000011000;
      15'b000_100001100101 : VALUE=19'b0000001_011000010111;
      15'b000_100001100110 : VALUE=19'b0000001_011000010110;
      15'b000_100001100111 : VALUE=19'b0000001_011000010100;
      15'b000_100001101000 : VALUE=19'b0000001_011000010011;
      15'b000_100001101001 : VALUE=19'b0000001_011000010010;
      15'b000_100001101010 : VALUE=19'b0000001_011000010000;
      15'b000_100001101011 : VALUE=19'b0000001_011000001111;
      15'b000_100001101100 : VALUE=19'b0000001_011000001110;
      15'b000_100001101101 : VALUE=19'b0000001_011000001100;
      15'b000_100001101110 : VALUE=19'b0000001_011000001011;
      15'b000_100001101111 : VALUE=19'b0000001_011000001010;
      15'b000_100001110000 : VALUE=19'b0000001_011000001000;
      15'b000_100001110001 : VALUE=19'b0000001_011000000111;
      15'b000_100001110010 : VALUE=19'b0000001_011000000110;
      15'b000_100001110011 : VALUE=19'b0000001_011000000101;
      15'b000_100001110100 : VALUE=19'b0000001_011000000011;
      15'b000_100001110101 : VALUE=19'b0000001_011000000010;
      15'b000_100001110110 : VALUE=19'b0000001_011000000001;
      15'b000_100001110111 : VALUE=19'b0000001_010111111111;
      15'b000_100001111000 : VALUE=19'b0000001_010111111110;
      15'b000_100001111001 : VALUE=19'b0000001_010111111101;
      15'b000_100001111010 : VALUE=19'b0000001_010111111011;
      15'b000_100001111011 : VALUE=19'b0000001_010111111010;
      15'b000_100001111100 : VALUE=19'b0000001_010111111001;
      15'b000_100001111101 : VALUE=19'b0000001_010111111000;
      15'b000_100001111110 : VALUE=19'b0000001_010111110110;
      15'b000_100001111111 : VALUE=19'b0000001_010111110101;
      15'b000_100010000000 : VALUE=19'b0000001_010111110100;
      15'b000_100010000001 : VALUE=19'b0000001_010111110010;
      15'b000_100010000010 : VALUE=19'b0000001_010111110001;
      15'b000_100010000011 : VALUE=19'b0000001_010111110000;
      15'b000_100010000100 : VALUE=19'b0000001_010111101111;
      15'b000_100010000101 : VALUE=19'b0000001_010111101101;
      15'b000_100010000110 : VALUE=19'b0000001_010111101100;
      15'b000_100010000111 : VALUE=19'b0000001_010111101011;
      15'b000_100010001000 : VALUE=19'b0000001_010111101001;
      15'b000_100010001001 : VALUE=19'b0000001_010111101000;
      15'b000_100010001010 : VALUE=19'b0000001_010111100111;
      15'b000_100010001011 : VALUE=19'b0000001_010111100110;
      15'b000_100010001100 : VALUE=19'b0000001_010111100100;
      15'b000_100010001101 : VALUE=19'b0000001_010111100011;
      15'b000_100010001110 : VALUE=19'b0000001_010111100010;
      15'b000_100010001111 : VALUE=19'b0000001_010111100000;
      15'b000_100010010000 : VALUE=19'b0000001_010111011111;
      15'b000_100010010001 : VALUE=19'b0000001_010111011110;
      15'b000_100010010010 : VALUE=19'b0000001_010111011101;
      15'b000_100010010011 : VALUE=19'b0000001_010111011011;
      15'b000_100010010100 : VALUE=19'b0000001_010111011010;
      15'b000_100010010101 : VALUE=19'b0000001_010111011001;
      15'b000_100010010110 : VALUE=19'b0000001_010111010111;
      15'b000_100010010111 : VALUE=19'b0000001_010111010110;
      15'b000_100010011000 : VALUE=19'b0000001_010111010101;
      15'b000_100010011001 : VALUE=19'b0000001_010111010100;
      15'b000_100010011010 : VALUE=19'b0000001_010111010010;
      15'b000_100010011011 : VALUE=19'b0000001_010111010001;
      15'b000_100010011100 : VALUE=19'b0000001_010111010000;
      15'b000_100010011101 : VALUE=19'b0000001_010111001111;
      15'b000_100010011110 : VALUE=19'b0000001_010111001101;
      15'b000_100010011111 : VALUE=19'b0000001_010111001100;
      15'b000_100010100000 : VALUE=19'b0000001_010111001011;
      15'b000_100010100001 : VALUE=19'b0000001_010111001010;
      15'b000_100010100010 : VALUE=19'b0000001_010111001000;
      15'b000_100010100011 : VALUE=19'b0000001_010111000111;
      15'b000_100010100100 : VALUE=19'b0000001_010111000110;
      15'b000_100010100101 : VALUE=19'b0000001_010111000100;
      15'b000_100010100110 : VALUE=19'b0000001_010111000011;
      15'b000_100010100111 : VALUE=19'b0000001_010111000010;
      15'b000_100010101000 : VALUE=19'b0000001_010111000001;
      15'b000_100010101001 : VALUE=19'b0000001_010110111111;
      15'b000_100010101010 : VALUE=19'b0000001_010110111110;
      15'b000_100010101011 : VALUE=19'b0000001_010110111101;
      15'b000_100010101100 : VALUE=19'b0000001_010110111100;
      15'b000_100010101101 : VALUE=19'b0000001_010110111010;
      15'b000_100010101110 : VALUE=19'b0000001_010110111001;
      15'b000_100010101111 : VALUE=19'b0000001_010110111000;
      15'b000_100010110000 : VALUE=19'b0000001_010110110111;
      15'b000_100010110001 : VALUE=19'b0000001_010110110101;
      15'b000_100010110010 : VALUE=19'b0000001_010110110100;
      15'b000_100010110011 : VALUE=19'b0000001_010110110011;
      15'b000_100010110100 : VALUE=19'b0000001_010110110010;
      15'b000_100010110101 : VALUE=19'b0000001_010110110000;
      15'b000_100010110110 : VALUE=19'b0000001_010110101111;
      15'b000_100010110111 : VALUE=19'b0000001_010110101110;
      15'b000_100010111000 : VALUE=19'b0000001_010110101101;
      15'b000_100010111001 : VALUE=19'b0000001_010110101011;
      15'b000_100010111010 : VALUE=19'b0000001_010110101010;
      15'b000_100010111011 : VALUE=19'b0000001_010110101001;
      15'b000_100010111100 : VALUE=19'b0000001_010110101000;
      15'b000_100010111101 : VALUE=19'b0000001_010110100111;
      15'b000_100010111110 : VALUE=19'b0000001_010110100101;
      15'b000_100010111111 : VALUE=19'b0000001_010110100100;
      15'b000_100011000000 : VALUE=19'b0000001_010110100011;
      15'b000_100011000001 : VALUE=19'b0000001_010110100010;
      15'b000_100011000010 : VALUE=19'b0000001_010110100000;
      15'b000_100011000011 : VALUE=19'b0000001_010110011111;
      15'b000_100011000100 : VALUE=19'b0000001_010110011110;
      15'b000_100011000101 : VALUE=19'b0000001_010110011101;
      15'b000_100011000110 : VALUE=19'b0000001_010110011011;
      15'b000_100011000111 : VALUE=19'b0000001_010110011010;
      15'b000_100011001000 : VALUE=19'b0000001_010110011001;
      15'b000_100011001001 : VALUE=19'b0000001_010110011000;
      15'b000_100011001010 : VALUE=19'b0000001_010110010110;
      15'b000_100011001011 : VALUE=19'b0000001_010110010101;
      15'b000_100011001100 : VALUE=19'b0000001_010110010100;
      15'b000_100011001101 : VALUE=19'b0000001_010110010011;
      15'b000_100011001110 : VALUE=19'b0000001_010110010010;
      15'b000_100011001111 : VALUE=19'b0000001_010110010000;
      15'b000_100011010000 : VALUE=19'b0000001_010110001111;
      15'b000_100011010001 : VALUE=19'b0000001_010110001110;
      15'b000_100011010010 : VALUE=19'b0000001_010110001101;
      15'b000_100011010011 : VALUE=19'b0000001_010110001011;
      15'b000_100011010100 : VALUE=19'b0000001_010110001010;
      15'b000_100011010101 : VALUE=19'b0000001_010110001001;
      15'b000_100011010110 : VALUE=19'b0000001_010110001000;
      15'b000_100011010111 : VALUE=19'b0000001_010110000111;
      15'b000_100011011000 : VALUE=19'b0000001_010110000101;
      15'b000_100011011001 : VALUE=19'b0000001_010110000100;
      15'b000_100011011010 : VALUE=19'b0000001_010110000011;
      15'b000_100011011011 : VALUE=19'b0000001_010110000010;
      15'b000_100011011100 : VALUE=19'b0000001_010110000001;
      15'b000_100011011101 : VALUE=19'b0000001_010101111111;
      15'b000_100011011110 : VALUE=19'b0000001_010101111110;
      15'b000_100011011111 : VALUE=19'b0000001_010101111101;
      15'b000_100011100000 : VALUE=19'b0000001_010101111100;
      15'b000_100011100001 : VALUE=19'b0000001_010101111010;
      15'b000_100011100010 : VALUE=19'b0000001_010101111001;
      15'b000_100011100011 : VALUE=19'b0000001_010101111000;
      15'b000_100011100100 : VALUE=19'b0000001_010101110111;
      15'b000_100011100101 : VALUE=19'b0000001_010101110110;
      15'b000_100011100110 : VALUE=19'b0000001_010101110100;
      15'b000_100011100111 : VALUE=19'b0000001_010101110011;
      15'b000_100011101000 : VALUE=19'b0000001_010101110010;
      15'b000_100011101001 : VALUE=19'b0000001_010101110001;
      15'b000_100011101010 : VALUE=19'b0000001_010101110000;
      15'b000_100011101011 : VALUE=19'b0000001_010101101110;
      15'b000_100011101100 : VALUE=19'b0000001_010101101101;
      15'b000_100011101101 : VALUE=19'b0000001_010101101100;
      15'b000_100011101110 : VALUE=19'b0000001_010101101011;
      15'b000_100011101111 : VALUE=19'b0000001_010101101010;
      15'b000_100011110000 : VALUE=19'b0000001_010101101000;
      15'b000_100011110001 : VALUE=19'b0000001_010101100111;
      15'b000_100011110010 : VALUE=19'b0000001_010101100110;
      15'b000_100011110011 : VALUE=19'b0000001_010101100101;
      15'b000_100011110100 : VALUE=19'b0000001_010101100100;
      15'b000_100011110101 : VALUE=19'b0000001_010101100010;
      15'b000_100011110110 : VALUE=19'b0000001_010101100001;
      15'b000_100011110111 : VALUE=19'b0000001_010101100000;
      15'b000_100011111000 : VALUE=19'b0000001_010101011111;
      15'b000_100011111001 : VALUE=19'b0000001_010101011110;
      15'b000_100011111010 : VALUE=19'b0000001_010101011100;
      15'b000_100011111011 : VALUE=19'b0000001_010101011011;
      15'b000_100011111100 : VALUE=19'b0000001_010101011010;
      15'b000_100011111101 : VALUE=19'b0000001_010101011001;
      15'b000_100011111110 : VALUE=19'b0000001_010101011000;
      15'b000_100011111111 : VALUE=19'b0000001_010101010111;
      15'b000_100100000000 : VALUE=19'b0000001_010101010101;
      15'b000_100100000001 : VALUE=19'b0000001_010101010100;
      15'b000_100100000010 : VALUE=19'b0000001_010101010011;
      15'b000_100100000011 : VALUE=19'b0000001_010101010010;
      15'b000_100100000100 : VALUE=19'b0000001_010101010001;
      15'b000_100100000101 : VALUE=19'b0000001_010101001111;
      15'b000_100100000110 : VALUE=19'b0000001_010101001110;
      15'b000_100100000111 : VALUE=19'b0000001_010101001101;
      15'b000_100100001000 : VALUE=19'b0000001_010101001100;
      15'b000_100100001001 : VALUE=19'b0000001_010101001011;
      15'b000_100100001010 : VALUE=19'b0000001_010101001010;
      15'b000_100100001011 : VALUE=19'b0000001_010101001000;
      15'b000_100100001100 : VALUE=19'b0000001_010101000111;
      15'b000_100100001101 : VALUE=19'b0000001_010101000110;
      15'b000_100100001110 : VALUE=19'b0000001_010101000101;
      15'b000_100100001111 : VALUE=19'b0000001_010101000100;
      15'b000_100100010000 : VALUE=19'b0000001_010101000010;
      15'b000_100100010001 : VALUE=19'b0000001_010101000001;
      15'b000_100100010010 : VALUE=19'b0000001_010101000000;
      15'b000_100100010011 : VALUE=19'b0000001_010100111111;
      15'b000_100100010100 : VALUE=19'b0000001_010100111110;
      15'b000_100100010101 : VALUE=19'b0000001_010100111101;
      15'b000_100100010110 : VALUE=19'b0000001_010100111011;
      15'b000_100100010111 : VALUE=19'b0000001_010100111010;
      15'b000_100100011000 : VALUE=19'b0000001_010100111001;
      15'b000_100100011001 : VALUE=19'b0000001_010100111000;
      15'b000_100100011010 : VALUE=19'b0000001_010100110111;
      15'b000_100100011011 : VALUE=19'b0000001_010100110110;
      15'b000_100100011100 : VALUE=19'b0000001_010100110100;
      15'b000_100100011101 : VALUE=19'b0000001_010100110011;
      15'b000_100100011110 : VALUE=19'b0000001_010100110010;
      15'b000_100100011111 : VALUE=19'b0000001_010100110001;
      15'b000_100100100000 : VALUE=19'b0000001_010100110000;
      15'b000_100100100001 : VALUE=19'b0000001_010100101111;
      15'b000_100100100010 : VALUE=19'b0000001_010100101101;
      15'b000_100100100011 : VALUE=19'b0000001_010100101100;
      15'b000_100100100100 : VALUE=19'b0000001_010100101011;
      15'b000_100100100101 : VALUE=19'b0000001_010100101010;
      15'b000_100100100110 : VALUE=19'b0000001_010100101001;
      15'b000_100100100111 : VALUE=19'b0000001_010100101000;
      15'b000_100100101000 : VALUE=19'b0000001_010100100111;
      15'b000_100100101001 : VALUE=19'b0000001_010100100101;
      15'b000_100100101010 : VALUE=19'b0000001_010100100100;
      15'b000_100100101011 : VALUE=19'b0000001_010100100011;
      15'b000_100100101100 : VALUE=19'b0000001_010100100010;
      15'b000_100100101101 : VALUE=19'b0000001_010100100001;
      15'b000_100100101110 : VALUE=19'b0000001_010100100000;
      15'b000_100100101111 : VALUE=19'b0000001_010100011110;
      15'b000_100100110000 : VALUE=19'b0000001_010100011101;
      15'b000_100100110001 : VALUE=19'b0000001_010100011100;
      15'b000_100100110010 : VALUE=19'b0000001_010100011011;
      15'b000_100100110011 : VALUE=19'b0000001_010100011010;
      15'b000_100100110100 : VALUE=19'b0000001_010100011001;
      15'b000_100100110101 : VALUE=19'b0000001_010100011000;
      15'b000_100100110110 : VALUE=19'b0000001_010100010110;
      15'b000_100100110111 : VALUE=19'b0000001_010100010101;
      15'b000_100100111000 : VALUE=19'b0000001_010100010100;
      15'b000_100100111001 : VALUE=19'b0000001_010100010011;
      15'b000_100100111010 : VALUE=19'b0000001_010100010010;
      15'b000_100100111011 : VALUE=19'b0000001_010100010001;
      15'b000_100100111100 : VALUE=19'b0000001_010100010000;
      15'b000_100100111101 : VALUE=19'b0000001_010100001110;
      15'b000_100100111110 : VALUE=19'b0000001_010100001101;
      15'b000_100100111111 : VALUE=19'b0000001_010100001100;
      15'b000_100101000000 : VALUE=19'b0000001_010100001011;
      15'b000_100101000001 : VALUE=19'b0000001_010100001010;
      15'b000_100101000010 : VALUE=19'b0000001_010100001001;
      15'b000_100101000011 : VALUE=19'b0000001_010100001000;
      15'b000_100101000100 : VALUE=19'b0000001_010100000110;
      15'b000_100101000101 : VALUE=19'b0000001_010100000101;
      15'b000_100101000110 : VALUE=19'b0000001_010100000100;
      15'b000_100101000111 : VALUE=19'b0000001_010100000011;
      15'b000_100101001000 : VALUE=19'b0000001_010100000010;
      15'b000_100101001001 : VALUE=19'b0000001_010100000001;
      15'b000_100101001010 : VALUE=19'b0000001_010100000000;
      15'b000_100101001011 : VALUE=19'b0000001_010011111111;
      15'b000_100101001100 : VALUE=19'b0000001_010011111101;
      15'b000_100101001101 : VALUE=19'b0000001_010011111100;
      15'b000_100101001110 : VALUE=19'b0000001_010011111011;
      15'b000_100101001111 : VALUE=19'b0000001_010011111010;
      15'b000_100101010000 : VALUE=19'b0000001_010011111001;
      15'b000_100101010001 : VALUE=19'b0000001_010011111000;
      15'b000_100101010010 : VALUE=19'b0000001_010011110111;
      15'b000_100101010011 : VALUE=19'b0000001_010011110110;
      15'b000_100101010100 : VALUE=19'b0000001_010011110100;
      15'b000_100101010101 : VALUE=19'b0000001_010011110011;
      15'b000_100101010110 : VALUE=19'b0000001_010011110010;
      15'b000_100101010111 : VALUE=19'b0000001_010011110001;
      15'b000_100101011000 : VALUE=19'b0000001_010011110000;
      15'b000_100101011001 : VALUE=19'b0000001_010011101111;
      15'b000_100101011010 : VALUE=19'b0000001_010011101110;
      15'b000_100101011011 : VALUE=19'b0000001_010011101101;
      15'b000_100101011100 : VALUE=19'b0000001_010011101011;
      15'b000_100101011101 : VALUE=19'b0000001_010011101010;
      15'b000_100101011110 : VALUE=19'b0000001_010011101001;
      15'b000_100101011111 : VALUE=19'b0000001_010011101000;
      15'b000_100101100000 : VALUE=19'b0000001_010011100111;
      15'b000_100101100001 : VALUE=19'b0000001_010011100110;
      15'b000_100101100010 : VALUE=19'b0000001_010011100101;
      15'b000_100101100011 : VALUE=19'b0000001_010011100100;
      15'b000_100101100100 : VALUE=19'b0000001_010011100011;
      15'b000_100101100101 : VALUE=19'b0000001_010011100001;
      15'b000_100101100110 : VALUE=19'b0000001_010011100000;
      15'b000_100101100111 : VALUE=19'b0000001_010011011111;
      15'b000_100101101000 : VALUE=19'b0000001_010011011110;
      15'b000_100101101001 : VALUE=19'b0000001_010011011101;
      15'b000_100101101010 : VALUE=19'b0000001_010011011100;
      15'b000_100101101011 : VALUE=19'b0000001_010011011011;
      15'b000_100101101100 : VALUE=19'b0000001_010011011010;
      15'b000_100101101101 : VALUE=19'b0000001_010011011001;
      15'b000_100101101110 : VALUE=19'b0000001_010011010111;
      15'b000_100101101111 : VALUE=19'b0000001_010011010110;
      15'b000_100101110000 : VALUE=19'b0000001_010011010101;
      15'b000_100101110001 : VALUE=19'b0000001_010011010100;
      15'b000_100101110010 : VALUE=19'b0000001_010011010011;
      15'b000_100101110011 : VALUE=19'b0000001_010011010010;
      15'b000_100101110100 : VALUE=19'b0000001_010011010001;
      15'b000_100101110101 : VALUE=19'b0000001_010011010000;
      15'b000_100101110110 : VALUE=19'b0000001_010011001111;
      15'b000_100101110111 : VALUE=19'b0000001_010011001110;
      15'b000_100101111000 : VALUE=19'b0000001_010011001100;
      15'b000_100101111001 : VALUE=19'b0000001_010011001011;
      15'b000_100101111010 : VALUE=19'b0000001_010011001010;
      15'b000_100101111011 : VALUE=19'b0000001_010011001001;
      15'b000_100101111100 : VALUE=19'b0000001_010011001000;
      15'b000_100101111101 : VALUE=19'b0000001_010011000111;
      15'b000_100101111110 : VALUE=19'b0000001_010011000110;
      15'b000_100101111111 : VALUE=19'b0000001_010011000101;
      15'b000_100110000000 : VALUE=19'b0000001_010011000100;
      15'b000_100110000001 : VALUE=19'b0000001_010011000011;
      15'b000_100110000010 : VALUE=19'b0000001_010011000001;
      15'b000_100110000011 : VALUE=19'b0000001_010011000000;
      15'b000_100110000100 : VALUE=19'b0000001_010010111111;
      15'b000_100110000101 : VALUE=19'b0000001_010010111110;
      15'b000_100110000110 : VALUE=19'b0000001_010010111101;
      15'b000_100110000111 : VALUE=19'b0000001_010010111100;
      15'b000_100110001000 : VALUE=19'b0000001_010010111011;
      15'b000_100110001001 : VALUE=19'b0000001_010010111010;
      15'b000_100110001010 : VALUE=19'b0000001_010010111001;
      15'b000_100110001011 : VALUE=19'b0000001_010010111000;
      15'b000_100110001100 : VALUE=19'b0000001_010010110111;
      15'b000_100110001101 : VALUE=19'b0000001_010010110110;
      15'b000_100110001110 : VALUE=19'b0000001_010010110100;
      15'b000_100110001111 : VALUE=19'b0000001_010010110011;
      15'b000_100110010000 : VALUE=19'b0000001_010010110010;
      15'b000_100110010001 : VALUE=19'b0000001_010010110001;
      15'b000_100110010010 : VALUE=19'b0000001_010010110000;
      15'b000_100110010011 : VALUE=19'b0000001_010010101111;
      15'b000_100110010100 : VALUE=19'b0000001_010010101110;
      15'b000_100110010101 : VALUE=19'b0000001_010010101101;
      15'b000_100110010110 : VALUE=19'b0000001_010010101100;
      15'b000_100110010111 : VALUE=19'b0000001_010010101011;
      15'b000_100110011000 : VALUE=19'b0000001_010010101010;
      15'b000_100110011001 : VALUE=19'b0000001_010010101001;
      15'b000_100110011010 : VALUE=19'b0000001_010010100111;
      15'b000_100110011011 : VALUE=19'b0000001_010010100110;
      15'b000_100110011100 : VALUE=19'b0000001_010010100101;
      15'b000_100110011101 : VALUE=19'b0000001_010010100100;
      15'b000_100110011110 : VALUE=19'b0000001_010010100011;
      15'b000_100110011111 : VALUE=19'b0000001_010010100010;
      15'b000_100110100000 : VALUE=19'b0000001_010010100001;
      15'b000_100110100001 : VALUE=19'b0000001_010010100000;
      15'b000_100110100010 : VALUE=19'b0000001_010010011111;
      15'b000_100110100011 : VALUE=19'b0000001_010010011110;
      15'b000_100110100100 : VALUE=19'b0000001_010010011101;
      15'b000_100110100101 : VALUE=19'b0000001_010010011100;
      15'b000_100110100110 : VALUE=19'b0000001_010010011011;
      15'b000_100110100111 : VALUE=19'b0000001_010010011010;
      15'b000_100110101000 : VALUE=19'b0000001_010010011000;
      15'b000_100110101001 : VALUE=19'b0000001_010010010111;
      15'b000_100110101010 : VALUE=19'b0000001_010010010110;
      15'b000_100110101011 : VALUE=19'b0000001_010010010101;
      15'b000_100110101100 : VALUE=19'b0000001_010010010100;
      15'b000_100110101101 : VALUE=19'b0000001_010010010011;
      15'b000_100110101110 : VALUE=19'b0000001_010010010010;
      15'b000_100110101111 : VALUE=19'b0000001_010010010001;
      15'b000_100110110000 : VALUE=19'b0000001_010010010000;
      15'b000_100110110001 : VALUE=19'b0000001_010010001111;
      15'b000_100110110010 : VALUE=19'b0000001_010010001110;
      15'b000_100110110011 : VALUE=19'b0000001_010010001101;
      15'b000_100110110100 : VALUE=19'b0000001_010010001100;
      15'b000_100110110101 : VALUE=19'b0000001_010010001011;
      15'b000_100110110110 : VALUE=19'b0000001_010010001010;
      15'b000_100110110111 : VALUE=19'b0000001_010010001001;
      15'b000_100110111000 : VALUE=19'b0000001_010010001000;
      15'b000_100110111001 : VALUE=19'b0000001_010010000110;
      15'b000_100110111010 : VALUE=19'b0000001_010010000101;
      15'b000_100110111011 : VALUE=19'b0000001_010010000100;
      15'b000_100110111100 : VALUE=19'b0000001_010010000011;
      15'b000_100110111101 : VALUE=19'b0000001_010010000010;
      15'b000_100110111110 : VALUE=19'b0000001_010010000001;
      15'b000_100110111111 : VALUE=19'b0000001_010010000000;
      15'b000_100111000000 : VALUE=19'b0000001_010001111111;
      15'b000_100111000001 : VALUE=19'b0000001_010001111110;
      15'b000_100111000010 : VALUE=19'b0000001_010001111101;
      15'b000_100111000011 : VALUE=19'b0000001_010001111100;
      15'b000_100111000100 : VALUE=19'b0000001_010001111011;
      15'b000_100111000101 : VALUE=19'b0000001_010001111010;
      15'b000_100111000110 : VALUE=19'b0000001_010001111001;
      15'b000_100111000111 : VALUE=19'b0000001_010001111000;
      15'b000_100111001000 : VALUE=19'b0000001_010001110111;
      15'b000_100111001001 : VALUE=19'b0000001_010001110110;
      15'b000_100111001010 : VALUE=19'b0000001_010001110101;
      15'b000_100111001011 : VALUE=19'b0000001_010001110100;
      15'b000_100111001100 : VALUE=19'b0000001_010001110011;
      15'b000_100111001101 : VALUE=19'b0000001_010001110001;
      15'b000_100111001110 : VALUE=19'b0000001_010001110000;
      15'b000_100111001111 : VALUE=19'b0000001_010001101111;
      15'b000_100111010000 : VALUE=19'b0000001_010001101110;
      15'b000_100111010001 : VALUE=19'b0000001_010001101101;
      15'b000_100111010010 : VALUE=19'b0000001_010001101100;
      15'b000_100111010011 : VALUE=19'b0000001_010001101011;
      15'b000_100111010100 : VALUE=19'b0000001_010001101010;
      15'b000_100111010101 : VALUE=19'b0000001_010001101001;
      15'b000_100111010110 : VALUE=19'b0000001_010001101000;
      15'b000_100111010111 : VALUE=19'b0000001_010001100111;
      15'b000_100111011000 : VALUE=19'b0000001_010001100110;
      15'b000_100111011001 : VALUE=19'b0000001_010001100101;
      15'b000_100111011010 : VALUE=19'b0000001_010001100100;
      15'b000_100111011011 : VALUE=19'b0000001_010001100011;
      15'b000_100111011100 : VALUE=19'b0000001_010001100010;
      15'b000_100111011101 : VALUE=19'b0000001_010001100001;
      15'b000_100111011110 : VALUE=19'b0000001_010001100000;
      15'b000_100111011111 : VALUE=19'b0000001_010001011111;
      15'b000_100111100000 : VALUE=19'b0000001_010001011110;
      15'b000_100111100001 : VALUE=19'b0000001_010001011101;
      15'b000_100111100010 : VALUE=19'b0000001_010001011100;
      15'b000_100111100011 : VALUE=19'b0000001_010001011011;
      15'b000_100111100100 : VALUE=19'b0000001_010001011010;
      15'b000_100111100101 : VALUE=19'b0000001_010001011001;
      15'b000_100111100110 : VALUE=19'b0000001_010001011000;
      15'b000_100111100111 : VALUE=19'b0000001_010001010111;
      15'b000_100111101000 : VALUE=19'b0000001_010001010110;
      15'b000_100111101001 : VALUE=19'b0000001_010001010101;
      15'b000_100111101010 : VALUE=19'b0000001_010001010011;
      15'b000_100111101011 : VALUE=19'b0000001_010001010010;
      15'b000_100111101100 : VALUE=19'b0000001_010001010001;
      15'b000_100111101101 : VALUE=19'b0000001_010001010000;
      15'b000_100111101110 : VALUE=19'b0000001_010001001111;
      15'b000_100111101111 : VALUE=19'b0000001_010001001110;
      15'b000_100111110000 : VALUE=19'b0000001_010001001101;
      15'b000_100111110001 : VALUE=19'b0000001_010001001100;
      15'b000_100111110010 : VALUE=19'b0000001_010001001011;
      15'b000_100111110011 : VALUE=19'b0000001_010001001010;
      15'b000_100111110100 : VALUE=19'b0000001_010001001001;
      15'b000_100111110101 : VALUE=19'b0000001_010001001000;
      15'b000_100111110110 : VALUE=19'b0000001_010001000111;
      15'b000_100111110111 : VALUE=19'b0000001_010001000110;
      15'b000_100111111000 : VALUE=19'b0000001_010001000101;
      15'b000_100111111001 : VALUE=19'b0000001_010001000100;
      15'b000_100111111010 : VALUE=19'b0000001_010001000011;
      15'b000_100111111011 : VALUE=19'b0000001_010001000010;
      15'b000_100111111100 : VALUE=19'b0000001_010001000001;
      15'b000_100111111101 : VALUE=19'b0000001_010001000000;
      15'b000_100111111110 : VALUE=19'b0000001_010000111111;
      15'b000_100111111111 : VALUE=19'b0000001_010000111110;
      15'b000_101000000000 : VALUE=19'b0000001_010000111101;
      15'b000_101000000001 : VALUE=19'b0000001_010000111100;
      15'b000_101000000010 : VALUE=19'b0000001_010000111011;
      15'b000_101000000011 : VALUE=19'b0000001_010000111010;
      15'b000_101000000100 : VALUE=19'b0000001_010000111001;
      15'b000_101000000101 : VALUE=19'b0000001_010000111000;
      15'b000_101000000110 : VALUE=19'b0000001_010000110111;
      15'b000_101000000111 : VALUE=19'b0000001_010000110110;
      15'b000_101000001000 : VALUE=19'b0000001_010000110101;
      15'b000_101000001001 : VALUE=19'b0000001_010000110100;
      15'b000_101000001010 : VALUE=19'b0000001_010000110011;
      15'b000_101000001011 : VALUE=19'b0000001_010000110010;
      15'b000_101000001100 : VALUE=19'b0000001_010000110001;
      15'b000_101000001101 : VALUE=19'b0000001_010000110000;
      15'b000_101000001110 : VALUE=19'b0000001_010000101111;
      15'b000_101000001111 : VALUE=19'b0000001_010000101110;
      15'b000_101000010000 : VALUE=19'b0000001_010000101101;
      15'b000_101000010001 : VALUE=19'b0000001_010000101100;
      15'b000_101000010010 : VALUE=19'b0000001_010000101011;
      15'b000_101000010011 : VALUE=19'b0000001_010000101010;
      15'b000_101000010100 : VALUE=19'b0000001_010000101001;
      15'b000_101000010101 : VALUE=19'b0000001_010000101000;
      15'b000_101000010110 : VALUE=19'b0000001_010000100111;
      15'b000_101000010111 : VALUE=19'b0000001_010000100110;
      15'b000_101000011000 : VALUE=19'b0000001_010000100101;
      15'b000_101000011001 : VALUE=19'b0000001_010000100100;
      15'b000_101000011010 : VALUE=19'b0000001_010000100011;
      15'b000_101000011011 : VALUE=19'b0000001_010000100010;
      15'b000_101000011100 : VALUE=19'b0000001_010000100001;
      15'b000_101000011101 : VALUE=19'b0000001_010000100000;
      15'b000_101000011110 : VALUE=19'b0000001_010000011111;
      15'b000_101000011111 : VALUE=19'b0000001_010000011110;
      15'b000_101000100000 : VALUE=19'b0000001_010000011101;
      15'b000_101000100001 : VALUE=19'b0000001_010000011100;
      15'b000_101000100010 : VALUE=19'b0000001_010000011011;
      15'b000_101000100011 : VALUE=19'b0000001_010000011010;
      15'b000_101000100100 : VALUE=19'b0000001_010000011001;
      15'b000_101000100101 : VALUE=19'b0000001_010000011000;
      15'b000_101000100110 : VALUE=19'b0000001_010000010111;
      15'b000_101000100111 : VALUE=19'b0000001_010000010110;
      15'b000_101000101000 : VALUE=19'b0000001_010000010101;
      15'b000_101000101001 : VALUE=19'b0000001_010000010100;
      15'b000_101000101010 : VALUE=19'b0000001_010000010011;
      15'b000_101000101011 : VALUE=19'b0000001_010000010010;
      15'b000_101000101100 : VALUE=19'b0000001_010000010001;
      15'b000_101000101101 : VALUE=19'b0000001_010000010000;
      15'b000_101000101110 : VALUE=19'b0000001_010000001111;
      15'b000_101000101111 : VALUE=19'b0000001_010000001110;
      15'b000_101000110000 : VALUE=19'b0000001_010000001101;
      15'b000_101000110001 : VALUE=19'b0000001_010000001100;
      15'b000_101000110010 : VALUE=19'b0000001_010000001011;
      15'b000_101000110011 : VALUE=19'b0000001_010000001010;
      15'b000_101000110100 : VALUE=19'b0000001_010000001001;
      15'b000_101000110101 : VALUE=19'b0000001_010000001000;
      15'b000_101000110110 : VALUE=19'b0000001_010000000111;
      15'b000_101000110111 : VALUE=19'b0000001_010000000110;
      15'b000_101000111000 : VALUE=19'b0000001_010000000101;
      15'b000_101000111001 : VALUE=19'b0000001_010000000100;
      15'b000_101000111010 : VALUE=19'b0000001_010000000011;
      15'b000_101000111011 : VALUE=19'b0000001_010000000010;
      15'b000_101000111100 : VALUE=19'b0000001_010000000001;
      15'b000_101000111101 : VALUE=19'b0000001_010000000000;
      15'b000_101000111110 : VALUE=19'b0000001_001111111111;
      15'b000_101000111111 : VALUE=19'b0000001_001111111110;
      15'b000_101001000000 : VALUE=19'b0000001_001111111110;
      15'b000_101001000001 : VALUE=19'b0000001_001111111101;
      15'b000_101001000010 : VALUE=19'b0000001_001111111100;
      15'b000_101001000011 : VALUE=19'b0000001_001111111011;
      15'b000_101001000100 : VALUE=19'b0000001_001111111010;
      15'b000_101001000101 : VALUE=19'b0000001_001111111001;
      15'b000_101001000110 : VALUE=19'b0000001_001111111000;
      15'b000_101001000111 : VALUE=19'b0000001_001111110111;
      15'b000_101001001000 : VALUE=19'b0000001_001111110110;
      15'b000_101001001001 : VALUE=19'b0000001_001111110101;
      15'b000_101001001010 : VALUE=19'b0000001_001111110100;
      15'b000_101001001011 : VALUE=19'b0000001_001111110011;
      15'b000_101001001100 : VALUE=19'b0000001_001111110010;
      15'b000_101001001101 : VALUE=19'b0000001_001111110001;
      15'b000_101001001110 : VALUE=19'b0000001_001111110000;
      15'b000_101001001111 : VALUE=19'b0000001_001111101111;
      15'b000_101001010000 : VALUE=19'b0000001_001111101110;
      15'b000_101001010001 : VALUE=19'b0000001_001111101101;
      15'b000_101001010010 : VALUE=19'b0000001_001111101100;
      15'b000_101001010011 : VALUE=19'b0000001_001111101011;
      15'b000_101001010100 : VALUE=19'b0000001_001111101010;
      15'b000_101001010101 : VALUE=19'b0000001_001111101001;
      15'b000_101001010110 : VALUE=19'b0000001_001111101000;
      15'b000_101001010111 : VALUE=19'b0000001_001111100111;
      15'b000_101001011000 : VALUE=19'b0000001_001111100110;
      15'b000_101001011001 : VALUE=19'b0000001_001111100101;
      15'b000_101001011010 : VALUE=19'b0000001_001111100100;
      15'b000_101001011011 : VALUE=19'b0000001_001111100011;
      15'b000_101001011100 : VALUE=19'b0000001_001111100010;
      15'b000_101001011101 : VALUE=19'b0000001_001111100001;
      15'b000_101001011110 : VALUE=19'b0000001_001111100000;
      15'b000_101001011111 : VALUE=19'b0000001_001111100000;
      15'b000_101001100000 : VALUE=19'b0000001_001111011111;
      15'b000_101001100001 : VALUE=19'b0000001_001111011110;
      15'b000_101001100010 : VALUE=19'b0000001_001111011101;
      15'b000_101001100011 : VALUE=19'b0000001_001111011100;
      15'b000_101001100100 : VALUE=19'b0000001_001111011011;
      15'b000_101001100101 : VALUE=19'b0000001_001111011010;
      15'b000_101001100110 : VALUE=19'b0000001_001111011001;
      15'b000_101001100111 : VALUE=19'b0000001_001111011000;
      15'b000_101001101000 : VALUE=19'b0000001_001111010111;
      15'b000_101001101001 : VALUE=19'b0000001_001111010110;
      15'b000_101001101010 : VALUE=19'b0000001_001111010101;
      15'b000_101001101011 : VALUE=19'b0000001_001111010100;
      15'b000_101001101100 : VALUE=19'b0000001_001111010011;
      15'b000_101001101101 : VALUE=19'b0000001_001111010010;
      15'b000_101001101110 : VALUE=19'b0000001_001111010001;
      15'b000_101001101111 : VALUE=19'b0000001_001111010000;
      15'b000_101001110000 : VALUE=19'b0000001_001111001111;
      15'b000_101001110001 : VALUE=19'b0000001_001111001110;
      15'b000_101001110010 : VALUE=19'b0000001_001111001101;
      15'b000_101001110011 : VALUE=19'b0000001_001111001100;
      15'b000_101001110100 : VALUE=19'b0000001_001111001100;
      15'b000_101001110101 : VALUE=19'b0000001_001111001011;
      15'b000_101001110110 : VALUE=19'b0000001_001111001010;
      15'b000_101001110111 : VALUE=19'b0000001_001111001001;
      15'b000_101001111000 : VALUE=19'b0000001_001111001000;
      15'b000_101001111001 : VALUE=19'b0000001_001111000111;
      15'b000_101001111010 : VALUE=19'b0000001_001111000110;
      15'b000_101001111011 : VALUE=19'b0000001_001111000101;
      15'b000_101001111100 : VALUE=19'b0000001_001111000100;
      15'b000_101001111101 : VALUE=19'b0000001_001111000011;
      15'b000_101001111110 : VALUE=19'b0000001_001111000010;
      15'b000_101001111111 : VALUE=19'b0000001_001111000001;
      15'b000_101010000000 : VALUE=19'b0000001_001111000000;
      15'b000_101010000001 : VALUE=19'b0000001_001110111111;
      15'b000_101010000010 : VALUE=19'b0000001_001110111110;
      15'b000_101010000011 : VALUE=19'b0000001_001110111101;
      15'b000_101010000100 : VALUE=19'b0000001_001110111100;
      15'b000_101010000101 : VALUE=19'b0000001_001110111100;
      15'b000_101010000110 : VALUE=19'b0000001_001110111011;
      15'b000_101010000111 : VALUE=19'b0000001_001110111010;
      15'b000_101010001000 : VALUE=19'b0000001_001110111001;
      15'b000_101010001001 : VALUE=19'b0000001_001110111000;
      15'b000_101010001010 : VALUE=19'b0000001_001110110111;
      15'b000_101010001011 : VALUE=19'b0000001_001110110110;
      15'b000_101010001100 : VALUE=19'b0000001_001110110101;
      15'b000_101010001101 : VALUE=19'b0000001_001110110100;
      15'b000_101010001110 : VALUE=19'b0000001_001110110011;
      15'b000_101010001111 : VALUE=19'b0000001_001110110010;
      15'b000_101010010000 : VALUE=19'b0000001_001110110001;
      15'b000_101010010001 : VALUE=19'b0000001_001110110000;
      15'b000_101010010010 : VALUE=19'b0000001_001110101111;
      15'b000_101010010011 : VALUE=19'b0000001_001110101110;
      15'b000_101010010100 : VALUE=19'b0000001_001110101110;
      15'b000_101010010101 : VALUE=19'b0000001_001110101101;
      15'b000_101010010110 : VALUE=19'b0000001_001110101100;
      15'b000_101010010111 : VALUE=19'b0000001_001110101011;
      15'b000_101010011000 : VALUE=19'b0000001_001110101010;
      15'b000_101010011001 : VALUE=19'b0000001_001110101001;
      15'b000_101010011010 : VALUE=19'b0000001_001110101000;
      15'b000_101010011011 : VALUE=19'b0000001_001110100111;
      15'b000_101010011100 : VALUE=19'b0000001_001110100110;
      15'b000_101010011101 : VALUE=19'b0000001_001110100101;
      15'b000_101010011110 : VALUE=19'b0000001_001110100100;
      15'b000_101010011111 : VALUE=19'b0000001_001110100011;
      15'b000_101010100000 : VALUE=19'b0000001_001110100010;
      15'b000_101010100001 : VALUE=19'b0000001_001110100001;
      15'b000_101010100010 : VALUE=19'b0000001_001110100001;
      15'b000_101010100011 : VALUE=19'b0000001_001110100000;
      15'b000_101010100100 : VALUE=19'b0000001_001110011111;
      15'b000_101010100101 : VALUE=19'b0000001_001110011110;
      15'b000_101010100110 : VALUE=19'b0000001_001110011101;
      15'b000_101010100111 : VALUE=19'b0000001_001110011100;
      15'b000_101010101000 : VALUE=19'b0000001_001110011011;
      15'b000_101010101001 : VALUE=19'b0000001_001110011010;
      15'b000_101010101010 : VALUE=19'b0000001_001110011001;
      15'b000_101010101011 : VALUE=19'b0000001_001110011000;
      15'b000_101010101100 : VALUE=19'b0000001_001110010111;
      15'b000_101010101101 : VALUE=19'b0000001_001110010110;
      15'b000_101010101110 : VALUE=19'b0000001_001110010101;
      15'b000_101010101111 : VALUE=19'b0000001_001110010101;
      15'b000_101010110000 : VALUE=19'b0000001_001110010100;
      15'b000_101010110001 : VALUE=19'b0000001_001110010011;
      15'b000_101010110010 : VALUE=19'b0000001_001110010010;
      15'b000_101010110011 : VALUE=19'b0000001_001110010001;
      15'b000_101010110100 : VALUE=19'b0000001_001110010000;
      15'b000_101010110101 : VALUE=19'b0000001_001110001111;
      15'b000_101010110110 : VALUE=19'b0000001_001110001110;
      15'b000_101010110111 : VALUE=19'b0000001_001110001101;
      15'b000_101010111000 : VALUE=19'b0000001_001110001100;
      15'b000_101010111001 : VALUE=19'b0000001_001110001011;
      15'b000_101010111010 : VALUE=19'b0000001_001110001011;
      15'b000_101010111011 : VALUE=19'b0000001_001110001010;
      15'b000_101010111100 : VALUE=19'b0000001_001110001001;
      15'b000_101010111101 : VALUE=19'b0000001_001110001000;
      15'b000_101010111110 : VALUE=19'b0000001_001110000111;
      15'b000_101010111111 : VALUE=19'b0000001_001110000110;
      15'b000_101011000000 : VALUE=19'b0000001_001110000101;
      15'b000_101011000001 : VALUE=19'b0000001_001110000100;
      15'b000_101011000010 : VALUE=19'b0000001_001110000011;
      15'b000_101011000011 : VALUE=19'b0000001_001110000010;
      15'b000_101011000100 : VALUE=19'b0000001_001110000001;
      15'b000_101011000101 : VALUE=19'b0000001_001110000001;
      15'b000_101011000110 : VALUE=19'b0000001_001110000000;
      15'b000_101011000111 : VALUE=19'b0000001_001101111111;
      15'b000_101011001000 : VALUE=19'b0000001_001101111110;
      15'b000_101011001001 : VALUE=19'b0000001_001101111101;
      15'b000_101011001010 : VALUE=19'b0000001_001101111100;
      15'b000_101011001011 : VALUE=19'b0000001_001101111011;
      15'b000_101011001100 : VALUE=19'b0000001_001101111010;
      15'b000_101011001101 : VALUE=19'b0000001_001101111001;
      15'b000_101011001110 : VALUE=19'b0000001_001101111000;
      15'b000_101011001111 : VALUE=19'b0000001_001101111000;
      15'b000_101011010000 : VALUE=19'b0000001_001101110111;
      15'b000_101011010001 : VALUE=19'b0000001_001101110110;
      15'b000_101011010010 : VALUE=19'b0000001_001101110101;
      15'b000_101011010011 : VALUE=19'b0000001_001101110100;
      15'b000_101011010100 : VALUE=19'b0000001_001101110011;
      15'b000_101011010101 : VALUE=19'b0000001_001101110010;
      15'b000_101011010110 : VALUE=19'b0000001_001101110001;
      15'b000_101011010111 : VALUE=19'b0000001_001101110000;
      15'b000_101011011000 : VALUE=19'b0000001_001101101111;
      15'b000_101011011001 : VALUE=19'b0000001_001101101111;
      15'b000_101011011010 : VALUE=19'b0000001_001101101110;
      15'b000_101011011011 : VALUE=19'b0000001_001101101101;
      15'b000_101011011100 : VALUE=19'b0000001_001101101100;
      15'b000_101011011101 : VALUE=19'b0000001_001101101011;
      15'b000_101011011110 : VALUE=19'b0000001_001101101010;
      15'b000_101011011111 : VALUE=19'b0000001_001101101001;
      15'b000_101011100000 : VALUE=19'b0000001_001101101000;
      15'b000_101011100001 : VALUE=19'b0000001_001101100111;
      15'b000_101011100010 : VALUE=19'b0000001_001101100110;
      15'b000_101011100011 : VALUE=19'b0000001_001101100110;
      15'b000_101011100100 : VALUE=19'b0000001_001101100101;
      15'b000_101011100101 : VALUE=19'b0000001_001101100100;
      15'b000_101011100110 : VALUE=19'b0000001_001101100011;
      15'b000_101011100111 : VALUE=19'b0000001_001101100010;
      15'b000_101011101000 : VALUE=19'b0000001_001101100001;
      15'b000_101011101001 : VALUE=19'b0000001_001101100000;
      15'b000_101011101010 : VALUE=19'b0000001_001101011111;
      15'b000_101011101011 : VALUE=19'b0000001_001101011110;
      15'b000_101011101100 : VALUE=19'b0000001_001101011110;
      15'b000_101011101101 : VALUE=19'b0000001_001101011101;
      15'b000_101011101110 : VALUE=19'b0000001_001101011100;
      15'b000_101011101111 : VALUE=19'b0000001_001101011011;
      15'b000_101011110000 : VALUE=19'b0000001_001101011010;
      15'b000_101011110001 : VALUE=19'b0000001_001101011001;
      15'b000_101011110010 : VALUE=19'b0000001_001101011000;
      15'b000_101011110011 : VALUE=19'b0000001_001101010111;
      15'b000_101011110100 : VALUE=19'b0000001_001101010111;
      15'b000_101011110101 : VALUE=19'b0000001_001101010110;
      15'b000_101011110110 : VALUE=19'b0000001_001101010101;
      15'b000_101011110111 : VALUE=19'b0000001_001101010100;
      15'b000_101011111000 : VALUE=19'b0000001_001101010011;
      15'b000_101011111001 : VALUE=19'b0000001_001101010010;
      15'b000_101011111010 : VALUE=19'b0000001_001101010001;
      15'b000_101011111011 : VALUE=19'b0000001_001101010000;
      15'b000_101011111100 : VALUE=19'b0000001_001101001111;
      15'b000_101011111101 : VALUE=19'b0000001_001101001111;
      15'b000_101011111110 : VALUE=19'b0000001_001101001110;
      15'b000_101011111111 : VALUE=19'b0000001_001101001101;
      15'b000_101100000000 : VALUE=19'b0000001_001101001100;
      15'b000_101100000001 : VALUE=19'b0000001_001101001011;
      15'b000_101100000010 : VALUE=19'b0000001_001101001010;
      15'b000_101100000011 : VALUE=19'b0000001_001101001001;
      15'b000_101100000100 : VALUE=19'b0000001_001101001000;
      15'b000_101100000101 : VALUE=19'b0000001_001101001000;
      15'b000_101100000110 : VALUE=19'b0000001_001101000111;
      15'b000_101100000111 : VALUE=19'b0000001_001101000110;
      15'b000_101100001000 : VALUE=19'b0000001_001101000101;
      15'b000_101100001001 : VALUE=19'b0000001_001101000100;
      15'b000_101100001010 : VALUE=19'b0000001_001101000011;
      15'b000_101100001011 : VALUE=19'b0000001_001101000010;
      15'b000_101100001100 : VALUE=19'b0000001_001101000001;
      15'b000_101100001101 : VALUE=19'b0000001_001101000001;
      15'b000_101100001110 : VALUE=19'b0000001_001101000000;
      15'b000_101100001111 : VALUE=19'b0000001_001100111111;
      15'b000_101100010000 : VALUE=19'b0000001_001100111110;
      15'b000_101100010001 : VALUE=19'b0000001_001100111101;
      15'b000_101100010010 : VALUE=19'b0000001_001100111100;
      15'b000_101100010011 : VALUE=19'b0000001_001100111011;
      15'b000_101100010100 : VALUE=19'b0000001_001100111011;
      15'b000_101100010101 : VALUE=19'b0000001_001100111010;
      15'b000_101100010110 : VALUE=19'b0000001_001100111001;
      15'b000_101100010111 : VALUE=19'b0000001_001100111000;
      15'b000_101100011000 : VALUE=19'b0000001_001100110111;
      15'b000_101100011001 : VALUE=19'b0000001_001100110110;
      15'b000_101100011010 : VALUE=19'b0000001_001100110101;
      15'b000_101100011011 : VALUE=19'b0000001_001100110100;
      15'b000_101100011100 : VALUE=19'b0000001_001100110100;
      15'b000_101100011101 : VALUE=19'b0000001_001100110011;
      15'b000_101100011110 : VALUE=19'b0000001_001100110010;
      15'b000_101100011111 : VALUE=19'b0000001_001100110001;
      15'b000_101100100000 : VALUE=19'b0000001_001100110000;
      15'b000_101100100001 : VALUE=19'b0000001_001100101111;
      15'b000_101100100010 : VALUE=19'b0000001_001100101110;
      15'b000_101100100011 : VALUE=19'b0000001_001100101110;
      15'b000_101100100100 : VALUE=19'b0000001_001100101101;
      15'b000_101100100101 : VALUE=19'b0000001_001100101100;
      15'b000_101100100110 : VALUE=19'b0000001_001100101011;
      15'b000_101100100111 : VALUE=19'b0000001_001100101010;
      15'b000_101100101000 : VALUE=19'b0000001_001100101001;
      15'b000_101100101001 : VALUE=19'b0000001_001100101000;
      15'b000_101100101010 : VALUE=19'b0000001_001100101000;
      15'b000_101100101011 : VALUE=19'b0000001_001100100111;
      15'b000_101100101100 : VALUE=19'b0000001_001100100110;
      15'b000_101100101101 : VALUE=19'b0000001_001100100101;
      15'b000_101100101110 : VALUE=19'b0000001_001100100100;
      15'b000_101100101111 : VALUE=19'b0000001_001100100011;
      15'b000_101100110000 : VALUE=19'b0000001_001100100010;
      15'b000_101100110001 : VALUE=19'b0000001_001100100010;
      15'b000_101100110010 : VALUE=19'b0000001_001100100001;
      15'b000_101100110011 : VALUE=19'b0000001_001100100000;
      15'b000_101100110100 : VALUE=19'b0000001_001100011111;
      15'b000_101100110101 : VALUE=19'b0000001_001100011110;
      15'b000_101100110110 : VALUE=19'b0000001_001100011101;
      15'b000_101100110111 : VALUE=19'b0000001_001100011100;
      15'b000_101100111000 : VALUE=19'b0000001_001100011100;
      15'b000_101100111001 : VALUE=19'b0000001_001100011011;
      15'b000_101100111010 : VALUE=19'b0000001_001100011010;
      15'b000_101100111011 : VALUE=19'b0000001_001100011001;
      15'b000_101100111100 : VALUE=19'b0000001_001100011000;
      15'b000_101100111101 : VALUE=19'b0000001_001100010111;
      15'b000_101100111110 : VALUE=19'b0000001_001100010110;
      15'b000_101100111111 : VALUE=19'b0000001_001100010110;
      15'b000_101101000000 : VALUE=19'b0000001_001100010101;
      15'b000_101101000001 : VALUE=19'b0000001_001100010100;
      15'b000_101101000010 : VALUE=19'b0000001_001100010011;
      15'b000_101101000011 : VALUE=19'b0000001_001100010010;
      15'b000_101101000100 : VALUE=19'b0000001_001100010001;
      15'b000_101101000101 : VALUE=19'b0000001_001100010001;
      15'b000_101101000110 : VALUE=19'b0000001_001100010000;
      15'b000_101101000111 : VALUE=19'b0000001_001100001111;
      15'b000_101101001000 : VALUE=19'b0000001_001100001110;
      15'b000_101101001001 : VALUE=19'b0000001_001100001101;
      15'b000_101101001010 : VALUE=19'b0000001_001100001100;
      15'b000_101101001011 : VALUE=19'b0000001_001100001011;
      15'b000_101101001100 : VALUE=19'b0000001_001100001011;
      15'b000_101101001101 : VALUE=19'b0000001_001100001010;
      15'b000_101101001110 : VALUE=19'b0000001_001100001001;
      15'b000_101101001111 : VALUE=19'b0000001_001100001000;
      15'b000_101101010000 : VALUE=19'b0000001_001100000111;
      15'b000_101101010001 : VALUE=19'b0000001_001100000110;
      15'b000_101101010010 : VALUE=19'b0000001_001100000110;
      15'b000_101101010011 : VALUE=19'b0000001_001100000101;
      15'b000_101101010100 : VALUE=19'b0000001_001100000100;
      15'b000_101101010101 : VALUE=19'b0000001_001100000011;
      15'b000_101101010110 : VALUE=19'b0000001_001100000010;
      15'b000_101101010111 : VALUE=19'b0000001_001100000001;
      15'b000_101101011000 : VALUE=19'b0000001_001100000001;
      15'b000_101101011001 : VALUE=19'b0000001_001100000000;
      15'b000_101101011010 : VALUE=19'b0000001_001011111111;
      15'b000_101101011011 : VALUE=19'b0000001_001011111110;
      15'b000_101101011100 : VALUE=19'b0000001_001011111101;
      15'b000_101101011101 : VALUE=19'b0000001_001011111100;
      15'b000_101101011110 : VALUE=19'b0000001_001011111100;
      15'b000_101101011111 : VALUE=19'b0000001_001011111011;
      15'b000_101101100000 : VALUE=19'b0000001_001011111010;
      15'b000_101101100001 : VALUE=19'b0000001_001011111001;
      15'b000_101101100010 : VALUE=19'b0000001_001011111000;
      15'b000_101101100011 : VALUE=19'b0000001_001011110111;
      15'b000_101101100100 : VALUE=19'b0000001_001011110111;
      15'b000_101101100101 : VALUE=19'b0000001_001011110110;
      15'b000_101101100110 : VALUE=19'b0000001_001011110101;
      15'b000_101101100111 : VALUE=19'b0000001_001011110100;
      15'b000_101101101000 : VALUE=19'b0000001_001011110011;
      15'b000_101101101001 : VALUE=19'b0000001_001011110010;
      15'b000_101101101010 : VALUE=19'b0000001_001011110010;
      15'b000_101101101011 : VALUE=19'b0000001_001011110001;
      15'b000_101101101100 : VALUE=19'b0000001_001011110000;
      15'b000_101101101101 : VALUE=19'b0000001_001011101111;
      15'b000_101101101110 : VALUE=19'b0000001_001011101110;
      15'b000_101101101111 : VALUE=19'b0000001_001011101101;
      15'b000_101101110000 : VALUE=19'b0000001_001011101101;
      15'b000_101101110001 : VALUE=19'b0000001_001011101100;
      15'b000_101101110010 : VALUE=19'b0000001_001011101011;
      15'b000_101101110011 : VALUE=19'b0000001_001011101010;
      15'b000_101101110100 : VALUE=19'b0000001_001011101001;
      15'b000_101101110101 : VALUE=19'b0000001_001011101000;
      15'b000_101101110110 : VALUE=19'b0000001_001011101000;
      15'b000_101101110111 : VALUE=19'b0000001_001011100111;
      15'b000_101101111000 : VALUE=19'b0000001_001011100110;
      15'b000_101101111001 : VALUE=19'b0000001_001011100101;
      15'b000_101101111010 : VALUE=19'b0000001_001011100100;
      15'b000_101101111011 : VALUE=19'b0000001_001011100011;
      15'b000_101101111100 : VALUE=19'b0000001_001011100011;
      15'b000_101101111101 : VALUE=19'b0000001_001011100010;
      15'b000_101101111110 : VALUE=19'b0000001_001011100001;
      15'b000_101101111111 : VALUE=19'b0000001_001011100000;
      15'b000_101110000000 : VALUE=19'b0000001_001011011111;
      15'b000_101110000001 : VALUE=19'b0000001_001011011111;
      15'b000_101110000010 : VALUE=19'b0000001_001011011110;
      15'b000_101110000011 : VALUE=19'b0000001_001011011101;
      15'b000_101110000100 : VALUE=19'b0000001_001011011100;
      15'b000_101110000101 : VALUE=19'b0000001_001011011011;
      15'b000_101110000110 : VALUE=19'b0000001_001011011010;
      15'b000_101110000111 : VALUE=19'b0000001_001011011010;
      15'b000_101110001000 : VALUE=19'b0000001_001011011001;
      15'b000_101110001001 : VALUE=19'b0000001_001011011000;
      15'b000_101110001010 : VALUE=19'b0000001_001011010111;
      15'b000_101110001011 : VALUE=19'b0000001_001011010110;
      15'b000_101110001100 : VALUE=19'b0000001_001011010110;
      15'b000_101110001101 : VALUE=19'b0000001_001011010101;
      15'b000_101110001110 : VALUE=19'b0000001_001011010100;
      15'b000_101110001111 : VALUE=19'b0000001_001011010011;
      15'b000_101110010000 : VALUE=19'b0000001_001011010010;
      15'b000_101110010001 : VALUE=19'b0000001_001011010001;
      15'b000_101110010010 : VALUE=19'b0000001_001011010001;
      15'b000_101110010011 : VALUE=19'b0000001_001011010000;
      15'b000_101110010100 : VALUE=19'b0000001_001011001111;
      15'b000_101110010101 : VALUE=19'b0000001_001011001110;
      15'b000_101110010110 : VALUE=19'b0000001_001011001101;
      15'b000_101110010111 : VALUE=19'b0000001_001011001101;
      15'b000_101110011000 : VALUE=19'b0000001_001011001100;
      15'b000_101110011001 : VALUE=19'b0000001_001011001011;
      15'b000_101110011010 : VALUE=19'b0000001_001011001010;
      15'b000_101110011011 : VALUE=19'b0000001_001011001001;
      15'b000_101110011100 : VALUE=19'b0000001_001011001001;
      15'b000_101110011101 : VALUE=19'b0000001_001011001000;
      15'b000_101110011110 : VALUE=19'b0000001_001011000111;
      15'b000_101110011111 : VALUE=19'b0000001_001011000110;
      15'b000_101110100000 : VALUE=19'b0000001_001011000101;
      15'b000_101110100001 : VALUE=19'b0000001_001011000101;
      15'b000_101110100010 : VALUE=19'b0000001_001011000100;
      15'b000_101110100011 : VALUE=19'b0000001_001011000011;
      15'b000_101110100100 : VALUE=19'b0000001_001011000010;
      15'b000_101110100101 : VALUE=19'b0000001_001011000001;
      15'b000_101110100110 : VALUE=19'b0000001_001011000000;
      15'b000_101110100111 : VALUE=19'b0000001_001011000000;
      15'b000_101110101000 : VALUE=19'b0000001_001010111111;
      15'b000_101110101001 : VALUE=19'b0000001_001010111110;
      15'b000_101110101010 : VALUE=19'b0000001_001010111101;
      15'b000_101110101011 : VALUE=19'b0000001_001010111100;
      15'b000_101110101100 : VALUE=19'b0000001_001010111100;
      15'b000_101110101101 : VALUE=19'b0000001_001010111011;
      15'b000_101110101110 : VALUE=19'b0000001_001010111010;
      15'b000_101110101111 : VALUE=19'b0000001_001010111001;
      15'b000_101110110000 : VALUE=19'b0000001_001010111000;
      15'b000_101110110001 : VALUE=19'b0000001_001010111000;
      15'b000_101110110010 : VALUE=19'b0000001_001010110111;
      15'b000_101110110011 : VALUE=19'b0000001_001010110110;
      15'b000_101110110100 : VALUE=19'b0000001_001010110101;
      15'b000_101110110101 : VALUE=19'b0000001_001010110100;
      15'b000_101110110110 : VALUE=19'b0000001_001010110100;
      15'b000_101110110111 : VALUE=19'b0000001_001010110011;
      15'b000_101110111000 : VALUE=19'b0000001_001010110010;
      15'b000_101110111001 : VALUE=19'b0000001_001010110001;
      15'b000_101110111010 : VALUE=19'b0000001_001010110000;
      15'b000_101110111011 : VALUE=19'b0000001_001010110000;
      15'b000_101110111100 : VALUE=19'b0000001_001010101111;
      15'b000_101110111101 : VALUE=19'b0000001_001010101110;
      15'b000_101110111110 : VALUE=19'b0000001_001010101101;
      15'b000_101110111111 : VALUE=19'b0000001_001010101100;
      15'b000_101111000000 : VALUE=19'b0000001_001010101100;
      15'b000_101111000001 : VALUE=19'b0000001_001010101011;
      15'b000_101111000010 : VALUE=19'b0000001_001010101010;
      15'b000_101111000011 : VALUE=19'b0000001_001010101001;
      15'b000_101111000100 : VALUE=19'b0000001_001010101001;
      15'b000_101111000101 : VALUE=19'b0000001_001010101000;
      15'b000_101111000110 : VALUE=19'b0000001_001010100111;
      15'b000_101111000111 : VALUE=19'b0000001_001010100110;
      15'b000_101111001000 : VALUE=19'b0000001_001010100101;
      15'b000_101111001001 : VALUE=19'b0000001_001010100101;
      15'b000_101111001010 : VALUE=19'b0000001_001010100100;
      15'b000_101111001011 : VALUE=19'b0000001_001010100011;
      15'b000_101111001100 : VALUE=19'b0000001_001010100010;
      15'b000_101111001101 : VALUE=19'b0000001_001010100001;
      15'b000_101111001110 : VALUE=19'b0000001_001010100001;
      15'b000_101111001111 : VALUE=19'b0000001_001010100000;
      15'b000_101111010000 : VALUE=19'b0000001_001010011111;
      15'b000_101111010001 : VALUE=19'b0000001_001010011110;
      15'b000_101111010010 : VALUE=19'b0000001_001010011101;
      15'b000_101111010011 : VALUE=19'b0000001_001010011101;
      15'b000_101111010100 : VALUE=19'b0000001_001010011100;
      15'b000_101111010101 : VALUE=19'b0000001_001010011011;
      15'b000_101111010110 : VALUE=19'b0000001_001010011010;
      15'b000_101111010111 : VALUE=19'b0000001_001010011010;
      15'b000_101111011000 : VALUE=19'b0000001_001010011001;
      15'b000_101111011001 : VALUE=19'b0000001_001010011000;
      15'b000_101111011010 : VALUE=19'b0000001_001010010111;
      15'b000_101111011011 : VALUE=19'b0000001_001010010110;
      15'b000_101111011100 : VALUE=19'b0000001_001010010110;
      15'b000_101111011101 : VALUE=19'b0000001_001010010101;
      15'b000_101111011110 : VALUE=19'b0000001_001010010100;
      15'b000_101111011111 : VALUE=19'b0000001_001010010011;
      15'b000_101111100000 : VALUE=19'b0000001_001010010010;
      15'b000_101111100001 : VALUE=19'b0000001_001010010010;
      15'b000_101111100010 : VALUE=19'b0000001_001010010001;
      15'b000_101111100011 : VALUE=19'b0000001_001010010000;
      15'b000_101111100100 : VALUE=19'b0000001_001010001111;
      15'b000_101111100101 : VALUE=19'b0000001_001010001111;
      15'b000_101111100110 : VALUE=19'b0000001_001010001110;
      15'b000_101111100111 : VALUE=19'b0000001_001010001101;
      15'b000_101111101000 : VALUE=19'b0000001_001010001100;
      15'b000_101111101001 : VALUE=19'b0000001_001010001011;
      15'b000_101111101010 : VALUE=19'b0000001_001010001011;
      15'b000_101111101011 : VALUE=19'b0000001_001010001010;
      15'b000_101111101100 : VALUE=19'b0000001_001010001001;
      15'b000_101111101101 : VALUE=19'b0000001_001010001000;
      15'b000_101111101110 : VALUE=19'b0000001_001010001000;
      15'b000_101111101111 : VALUE=19'b0000001_001010000111;
      15'b000_101111110000 : VALUE=19'b0000001_001010000110;
      15'b000_101111110001 : VALUE=19'b0000001_001010000101;
      15'b000_101111110010 : VALUE=19'b0000001_001010000100;
      15'b000_101111110011 : VALUE=19'b0000001_001010000100;
      15'b000_101111110100 : VALUE=19'b0000001_001010000011;
      15'b000_101111110101 : VALUE=19'b0000001_001010000010;
      15'b000_101111110110 : VALUE=19'b0000001_001010000001;
      15'b000_101111110111 : VALUE=19'b0000001_001010000001;
      15'b000_101111111000 : VALUE=19'b0000001_001010000000;
      15'b000_101111111001 : VALUE=19'b0000001_001001111111;
      15'b000_101111111010 : VALUE=19'b0000001_001001111110;
      15'b000_101111111011 : VALUE=19'b0000001_001001111110;
      15'b000_101111111100 : VALUE=19'b0000001_001001111101;
      15'b000_101111111101 : VALUE=19'b0000001_001001111100;
      15'b000_101111111110 : VALUE=19'b0000001_001001111011;
      15'b000_101111111111 : VALUE=19'b0000001_001001111010;
      15'b000_110000000000 : VALUE=19'b0000001_001001111010;
      15'b000_110000000001 : VALUE=19'b0000001_001001111001;
      15'b000_110000000010 : VALUE=19'b0000001_001001111000;
      15'b000_110000000011 : VALUE=19'b0000001_001001110111;
      15'b000_110000000100 : VALUE=19'b0000001_001001110111;
      15'b000_110000000101 : VALUE=19'b0000001_001001110110;
      15'b000_110000000110 : VALUE=19'b0000001_001001110101;
      15'b000_110000000111 : VALUE=19'b0000001_001001110100;
      15'b000_110000001000 : VALUE=19'b0000001_001001110100;
      15'b000_110000001001 : VALUE=19'b0000001_001001110011;
      15'b000_110000001010 : VALUE=19'b0000001_001001110010;
      15'b000_110000001011 : VALUE=19'b0000001_001001110001;
      15'b000_110000001100 : VALUE=19'b0000001_001001110000;
      15'b000_110000001101 : VALUE=19'b0000001_001001110000;
      15'b000_110000001110 : VALUE=19'b0000001_001001101111;
      15'b000_110000001111 : VALUE=19'b0000001_001001101110;
      15'b000_110000010000 : VALUE=19'b0000001_001001101101;
      15'b000_110000010001 : VALUE=19'b0000001_001001101101;
      15'b000_110000010010 : VALUE=19'b0000001_001001101100;
      15'b000_110000010011 : VALUE=19'b0000001_001001101011;
      15'b000_110000010100 : VALUE=19'b0000001_001001101010;
      15'b000_110000010101 : VALUE=19'b0000001_001001101010;
      15'b000_110000010110 : VALUE=19'b0000001_001001101001;
      15'b000_110000010111 : VALUE=19'b0000001_001001101000;
      15'b000_110000011000 : VALUE=19'b0000001_001001100111;
      15'b000_110000011001 : VALUE=19'b0000001_001001100111;
      15'b000_110000011010 : VALUE=19'b0000001_001001100110;
      15'b000_110000011011 : VALUE=19'b0000001_001001100101;
      15'b000_110000011100 : VALUE=19'b0000001_001001100100;
      15'b000_110000011101 : VALUE=19'b0000001_001001100011;
      15'b000_110000011110 : VALUE=19'b0000001_001001100011;
      15'b000_110000011111 : VALUE=19'b0000001_001001100010;
      15'b000_110000100000 : VALUE=19'b0000001_001001100001;
      15'b000_110000100001 : VALUE=19'b0000001_001001100000;
      15'b000_110000100010 : VALUE=19'b0000001_001001100000;
      15'b000_110000100011 : VALUE=19'b0000001_001001011111;
      15'b000_110000100100 : VALUE=19'b0000001_001001011110;
      15'b000_110000100101 : VALUE=19'b0000001_001001011101;
      15'b000_110000100110 : VALUE=19'b0000001_001001011101;
      15'b000_110000100111 : VALUE=19'b0000001_001001011100;
      15'b000_110000101000 : VALUE=19'b0000001_001001011011;
      15'b000_110000101001 : VALUE=19'b0000001_001001011010;
      15'b000_110000101010 : VALUE=19'b0000001_001001011010;
      15'b000_110000101011 : VALUE=19'b0000001_001001011001;
      15'b000_110000101100 : VALUE=19'b0000001_001001011000;
      15'b000_110000101101 : VALUE=19'b0000001_001001010111;
      15'b000_110000101110 : VALUE=19'b0000001_001001010111;
      15'b000_110000101111 : VALUE=19'b0000001_001001010110;
      15'b000_110000110000 : VALUE=19'b0000001_001001010101;
      15'b000_110000110001 : VALUE=19'b0000001_001001010100;
      15'b000_110000110010 : VALUE=19'b0000001_001001010100;
      15'b000_110000110011 : VALUE=19'b0000001_001001010011;
      15'b000_110000110100 : VALUE=19'b0000001_001001010010;
      15'b000_110000110101 : VALUE=19'b0000001_001001010001;
      15'b000_110000110110 : VALUE=19'b0000001_001001010001;
      15'b000_110000110111 : VALUE=19'b0000001_001001010000;
      15'b000_110000111000 : VALUE=19'b0000001_001001001111;
      15'b000_110000111001 : VALUE=19'b0000001_001001001110;
      15'b000_110000111010 : VALUE=19'b0000001_001001001110;
      15'b000_110000111011 : VALUE=19'b0000001_001001001101;
      15'b000_110000111100 : VALUE=19'b0000001_001001001100;
      15'b000_110000111101 : VALUE=19'b0000001_001001001011;
      15'b000_110000111110 : VALUE=19'b0000001_001001001011;
      15'b000_110000111111 : VALUE=19'b0000001_001001001010;
      15'b000_110001000000 : VALUE=19'b0000001_001001001001;
      15'b000_110001000001 : VALUE=19'b0000001_001001001000;
      15'b000_110001000010 : VALUE=19'b0000001_001001001000;
      15'b000_110001000011 : VALUE=19'b0000001_001001000111;
      15'b000_110001000100 : VALUE=19'b0000001_001001000110;
      15'b000_110001000101 : VALUE=19'b0000001_001001000101;
      15'b000_110001000110 : VALUE=19'b0000001_001001000101;
      15'b000_110001000111 : VALUE=19'b0000001_001001000100;
      15'b000_110001001000 : VALUE=19'b0000001_001001000011;
      15'b000_110001001001 : VALUE=19'b0000001_001001000010;
      15'b000_110001001010 : VALUE=19'b0000001_001001000010;
      15'b000_110001001011 : VALUE=19'b0000001_001001000001;
      15'b000_110001001100 : VALUE=19'b0000001_001001000000;
      15'b000_110001001101 : VALUE=19'b0000001_001000111111;
      15'b000_110001001110 : VALUE=19'b0000001_001000111111;
      15'b000_110001001111 : VALUE=19'b0000001_001000111110;
      15'b000_110001010000 : VALUE=19'b0000001_001000111101;
      15'b000_110001010001 : VALUE=19'b0000001_001000111101;
      15'b000_110001010010 : VALUE=19'b0000001_001000111100;
      15'b000_110001010011 : VALUE=19'b0000001_001000111011;
      15'b000_110001010100 : VALUE=19'b0000001_001000111010;
      15'b000_110001010101 : VALUE=19'b0000001_001000111010;
      15'b000_110001010110 : VALUE=19'b0000001_001000111001;
      15'b000_110001010111 : VALUE=19'b0000001_001000111000;
      15'b000_110001011000 : VALUE=19'b0000001_001000110111;
      15'b000_110001011001 : VALUE=19'b0000001_001000110111;
      15'b000_110001011010 : VALUE=19'b0000001_001000110110;
      15'b000_110001011011 : VALUE=19'b0000001_001000110101;
      15'b000_110001011100 : VALUE=19'b0000001_001000110100;
      15'b000_110001011101 : VALUE=19'b0000001_001000110100;
      15'b000_110001011110 : VALUE=19'b0000001_001000110011;
      15'b000_110001011111 : VALUE=19'b0000001_001000110010;
      15'b000_110001100000 : VALUE=19'b0000001_001000110001;
      15'b000_110001100001 : VALUE=19'b0000001_001000110001;
      15'b000_110001100010 : VALUE=19'b0000001_001000110000;
      15'b000_110001100011 : VALUE=19'b0000001_001000101111;
      15'b000_110001100100 : VALUE=19'b0000001_001000101111;
      15'b000_110001100101 : VALUE=19'b0000001_001000101110;
      15'b000_110001100110 : VALUE=19'b0000001_001000101101;
      15'b000_110001100111 : VALUE=19'b0000001_001000101100;
      15'b000_110001101000 : VALUE=19'b0000001_001000101100;
      15'b000_110001101001 : VALUE=19'b0000001_001000101011;
      15'b000_110001101010 : VALUE=19'b0000001_001000101010;
      15'b000_110001101011 : VALUE=19'b0000001_001000101001;
      15'b000_110001101100 : VALUE=19'b0000001_001000101001;
      15'b000_110001101101 : VALUE=19'b0000001_001000101000;
      15'b000_110001101110 : VALUE=19'b0000001_001000100111;
      15'b000_110001101111 : VALUE=19'b0000001_001000100110;
      15'b000_110001110000 : VALUE=19'b0000001_001000100110;
      15'b000_110001110001 : VALUE=19'b0000001_001000100101;
      15'b000_110001110010 : VALUE=19'b0000001_001000100100;
      15'b000_110001110011 : VALUE=19'b0000001_001000100100;
      15'b000_110001110100 : VALUE=19'b0000001_001000100011;
      15'b000_110001110101 : VALUE=19'b0000001_001000100010;
      15'b000_110001110110 : VALUE=19'b0000001_001000100001;
      15'b000_110001110111 : VALUE=19'b0000001_001000100001;
      15'b000_110001111000 : VALUE=19'b0000001_001000100000;
      15'b000_110001111001 : VALUE=19'b0000001_001000011111;
      15'b000_110001111010 : VALUE=19'b0000001_001000011110;
      15'b000_110001111011 : VALUE=19'b0000001_001000011110;
      15'b000_110001111100 : VALUE=19'b0000001_001000011101;
      15'b000_110001111101 : VALUE=19'b0000001_001000011100;
      15'b000_110001111110 : VALUE=19'b0000001_001000011100;
      15'b000_110001111111 : VALUE=19'b0000001_001000011011;
      15'b000_110010000000 : VALUE=19'b0000001_001000011010;
      15'b000_110010000001 : VALUE=19'b0000001_001000011001;
      15'b000_110010000010 : VALUE=19'b0000001_001000011001;
      15'b000_110010000011 : VALUE=19'b0000001_001000011000;
      15'b000_110010000100 : VALUE=19'b0000001_001000010111;
      15'b000_110010000101 : VALUE=19'b0000001_001000010110;
      15'b000_110010000110 : VALUE=19'b0000001_001000010110;
      15'b000_110010000111 : VALUE=19'b0000001_001000010101;
      15'b000_110010001000 : VALUE=19'b0000001_001000010100;
      15'b000_110010001001 : VALUE=19'b0000001_001000010100;
      15'b000_110010001010 : VALUE=19'b0000001_001000010011;
      15'b000_110010001011 : VALUE=19'b0000001_001000010010;
      15'b000_110010001100 : VALUE=19'b0000001_001000010001;
      15'b000_110010001101 : VALUE=19'b0000001_001000010001;
      15'b000_110010001110 : VALUE=19'b0000001_001000010000;
      15'b000_110010001111 : VALUE=19'b0000001_001000001111;
      15'b000_110010010000 : VALUE=19'b0000001_001000001111;
      15'b000_110010010001 : VALUE=19'b0000001_001000001110;
      15'b000_110010010010 : VALUE=19'b0000001_001000001101;
      15'b000_110010010011 : VALUE=19'b0000001_001000001100;
      15'b000_110010010100 : VALUE=19'b0000001_001000001100;
      15'b000_110010010101 : VALUE=19'b0000001_001000001011;
      15'b000_110010010110 : VALUE=19'b0000001_001000001010;
      15'b000_110010010111 : VALUE=19'b0000001_001000001010;
      15'b000_110010011000 : VALUE=19'b0000001_001000001001;
      15'b000_110010011001 : VALUE=19'b0000001_001000001000;
      15'b000_110010011010 : VALUE=19'b0000001_001000000111;
      15'b000_110010011011 : VALUE=19'b0000001_001000000111;
      15'b000_110010011100 : VALUE=19'b0000001_001000000110;
      15'b000_110010011101 : VALUE=19'b0000001_001000000101;
      15'b000_110010011110 : VALUE=19'b0000001_001000000101;
      15'b000_110010011111 : VALUE=19'b0000001_001000000100;
      15'b000_110010100000 : VALUE=19'b0000001_001000000011;
      15'b000_110010100001 : VALUE=19'b0000001_001000000010;
      15'b000_110010100010 : VALUE=19'b0000001_001000000010;
      15'b000_110010100011 : VALUE=19'b0000001_001000000001;
      15'b000_110010100100 : VALUE=19'b0000001_001000000000;
      15'b000_110010100101 : VALUE=19'b0000001_001000000000;
      15'b000_110010100110 : VALUE=19'b0000001_000111111111;
      15'b000_110010100111 : VALUE=19'b0000001_000111111110;
      15'b000_110010101000 : VALUE=19'b0000001_000111111101;
      15'b000_110010101001 : VALUE=19'b0000001_000111111101;
      15'b000_110010101010 : VALUE=19'b0000001_000111111100;
      15'b000_110010101011 : VALUE=19'b0000001_000111111011;
      15'b000_110010101100 : VALUE=19'b0000001_000111111011;
      15'b000_110010101101 : VALUE=19'b0000001_000111111010;
      15'b000_110010101110 : VALUE=19'b0000001_000111111001;
      15'b000_110010101111 : VALUE=19'b0000001_000111111000;
      15'b000_110010110000 : VALUE=19'b0000001_000111111000;
      15'b000_110010110001 : VALUE=19'b0000001_000111110111;
      15'b000_110010110010 : VALUE=19'b0000001_000111110110;
      15'b000_110010110011 : VALUE=19'b0000001_000111110110;
      15'b000_110010110100 : VALUE=19'b0000001_000111110101;
      15'b000_110010110101 : VALUE=19'b0000001_000111110100;
      15'b000_110010110110 : VALUE=19'b0000001_000111110011;
      15'b000_110010110111 : VALUE=19'b0000001_000111110011;
      15'b000_110010111000 : VALUE=19'b0000001_000111110010;
      15'b000_110010111001 : VALUE=19'b0000001_000111110001;
      15'b000_110010111010 : VALUE=19'b0000001_000111110001;
      15'b000_110010111011 : VALUE=19'b0000001_000111110000;
      15'b000_110010111100 : VALUE=19'b0000001_000111101111;
      15'b000_110010111101 : VALUE=19'b0000001_000111101111;
      15'b000_110010111110 : VALUE=19'b0000001_000111101110;
      15'b000_110010111111 : VALUE=19'b0000001_000111101101;
      15'b000_110011000000 : VALUE=19'b0000001_000111101100;
      15'b000_110011000001 : VALUE=19'b0000001_000111101100;
      15'b000_110011000010 : VALUE=19'b0000001_000111101011;
      15'b000_110011000011 : VALUE=19'b0000001_000111101010;
      15'b000_110011000100 : VALUE=19'b0000001_000111101010;
      15'b000_110011000101 : VALUE=19'b0000001_000111101001;
      15'b000_110011000110 : VALUE=19'b0000001_000111101000;
      15'b000_110011000111 : VALUE=19'b0000001_000111101000;
      15'b000_110011001000 : VALUE=19'b0000001_000111100111;
      15'b000_110011001001 : VALUE=19'b0000001_000111100110;
      15'b000_110011001010 : VALUE=19'b0000001_000111100101;
      15'b000_110011001011 : VALUE=19'b0000001_000111100101;
      15'b000_110011001100 : VALUE=19'b0000001_000111100100;
      15'b000_110011001101 : VALUE=19'b0000001_000111100011;
      15'b000_110011001110 : VALUE=19'b0000001_000111100011;
      15'b000_110011001111 : VALUE=19'b0000001_000111100010;
      15'b000_110011010000 : VALUE=19'b0000001_000111100001;
      15'b000_110011010001 : VALUE=19'b0000001_000111100001;
      15'b000_110011010010 : VALUE=19'b0000001_000111100000;
      15'b000_110011010011 : VALUE=19'b0000001_000111011111;
      15'b000_110011010100 : VALUE=19'b0000001_000111011110;
      15'b000_110011010101 : VALUE=19'b0000001_000111011110;
      15'b000_110011010110 : VALUE=19'b0000001_000111011101;
      15'b000_110011010111 : VALUE=19'b0000001_000111011100;
      15'b000_110011011000 : VALUE=19'b0000001_000111011100;
      15'b000_110011011001 : VALUE=19'b0000001_000111011011;
      15'b000_110011011010 : VALUE=19'b0000001_000111011010;
      15'b000_110011011011 : VALUE=19'b0000001_000111011010;
      15'b000_110011011100 : VALUE=19'b0000001_000111011001;
      15'b000_110011011101 : VALUE=19'b0000001_000111011000;
      15'b000_110011011110 : VALUE=19'b0000001_000111010111;
      15'b000_110011011111 : VALUE=19'b0000001_000111010111;
      15'b000_110011100000 : VALUE=19'b0000001_000111010110;
      15'b000_110011100001 : VALUE=19'b0000001_000111010101;
      15'b000_110011100010 : VALUE=19'b0000001_000111010101;
      15'b000_110011100011 : VALUE=19'b0000001_000111010100;
      15'b000_110011100100 : VALUE=19'b0000001_000111010011;
      15'b000_110011100101 : VALUE=19'b0000001_000111010011;
      15'b000_110011100110 : VALUE=19'b0000001_000111010010;
      15'b000_110011100111 : VALUE=19'b0000001_000111010001;
      15'b000_110011101000 : VALUE=19'b0000001_000111010001;
      15'b000_110011101001 : VALUE=19'b0000001_000111010000;
      15'b000_110011101010 : VALUE=19'b0000001_000111001111;
      15'b000_110011101011 : VALUE=19'b0000001_000111001111;
      15'b000_110011101100 : VALUE=19'b0000001_000111001110;
      15'b000_110011101101 : VALUE=19'b0000001_000111001101;
      15'b000_110011101110 : VALUE=19'b0000001_000111001100;
      15'b000_110011101111 : VALUE=19'b0000001_000111001100;
      15'b000_110011110000 : VALUE=19'b0000001_000111001011;
      15'b000_110011110001 : VALUE=19'b0000001_000111001010;
      15'b000_110011110010 : VALUE=19'b0000001_000111001010;
      15'b000_110011110011 : VALUE=19'b0000001_000111001001;
      15'b000_110011110100 : VALUE=19'b0000001_000111001000;
      15'b000_110011110101 : VALUE=19'b0000001_000111001000;
      15'b000_110011110110 : VALUE=19'b0000001_000111000111;
      15'b000_110011110111 : VALUE=19'b0000001_000111000110;
      15'b000_110011111000 : VALUE=19'b0000001_000111000110;
      15'b000_110011111001 : VALUE=19'b0000001_000111000101;
      15'b000_110011111010 : VALUE=19'b0000001_000111000100;
      15'b000_110011111011 : VALUE=19'b0000001_000111000100;
      15'b000_110011111100 : VALUE=19'b0000001_000111000011;
      15'b000_110011111101 : VALUE=19'b0000001_000111000010;
      15'b000_110011111110 : VALUE=19'b0000001_000111000001;
      15'b000_110011111111 : VALUE=19'b0000001_000111000001;
      15'b000_110100000000 : VALUE=19'b0000001_000111000000;
      15'b000_110100000001 : VALUE=19'b0000001_000110111111;
      15'b000_110100000010 : VALUE=19'b0000001_000110111111;
      15'b000_110100000011 : VALUE=19'b0000001_000110111110;
      15'b000_110100000100 : VALUE=19'b0000001_000110111101;
      15'b000_110100000101 : VALUE=19'b0000001_000110111101;
      15'b000_110100000110 : VALUE=19'b0000001_000110111100;
      15'b000_110100000111 : VALUE=19'b0000001_000110111011;
      15'b000_110100001000 : VALUE=19'b0000001_000110111011;
      15'b000_110100001001 : VALUE=19'b0000001_000110111010;
      15'b000_110100001010 : VALUE=19'b0000001_000110111001;
      15'b000_110100001011 : VALUE=19'b0000001_000110111001;
      15'b000_110100001100 : VALUE=19'b0000001_000110111000;
      15'b000_110100001101 : VALUE=19'b0000001_000110110111;
      15'b000_110100001110 : VALUE=19'b0000001_000110110111;
      15'b000_110100001111 : VALUE=19'b0000001_000110110110;
      15'b000_110100010000 : VALUE=19'b0000001_000110110101;
      15'b000_110100010001 : VALUE=19'b0000001_000110110101;
      15'b000_110100010010 : VALUE=19'b0000001_000110110100;
      15'b000_110100010011 : VALUE=19'b0000001_000110110011;
      15'b000_110100010100 : VALUE=19'b0000001_000110110011;
      15'b000_110100010101 : VALUE=19'b0000001_000110110010;
      15'b000_110100010110 : VALUE=19'b0000001_000110110001;
      15'b000_110100010111 : VALUE=19'b0000001_000110110000;
      15'b000_110100011000 : VALUE=19'b0000001_000110110000;
      15'b000_110100011001 : VALUE=19'b0000001_000110101111;
      15'b000_110100011010 : VALUE=19'b0000001_000110101110;
      15'b000_110100011011 : VALUE=19'b0000001_000110101110;
      15'b000_110100011100 : VALUE=19'b0000001_000110101101;
      15'b000_110100011101 : VALUE=19'b0000001_000110101100;
      15'b000_110100011110 : VALUE=19'b0000001_000110101100;
      15'b000_110100011111 : VALUE=19'b0000001_000110101011;
      15'b000_110100100000 : VALUE=19'b0000001_000110101010;
      15'b000_110100100001 : VALUE=19'b0000001_000110101010;
      15'b000_110100100010 : VALUE=19'b0000001_000110101001;
      15'b000_110100100011 : VALUE=19'b0000001_000110101000;
      15'b000_110100100100 : VALUE=19'b0000001_000110101000;
      15'b000_110100100101 : VALUE=19'b0000001_000110100111;
      15'b000_110100100110 : VALUE=19'b0000001_000110100110;
      15'b000_110100100111 : VALUE=19'b0000001_000110100110;
      15'b000_110100101000 : VALUE=19'b0000001_000110100101;
      15'b000_110100101001 : VALUE=19'b0000001_000110100100;
      15'b000_110100101010 : VALUE=19'b0000001_000110100100;
      15'b000_110100101011 : VALUE=19'b0000001_000110100011;
      15'b000_110100101100 : VALUE=19'b0000001_000110100010;
      15'b000_110100101101 : VALUE=19'b0000001_000110100010;
      15'b000_110100101110 : VALUE=19'b0000001_000110100001;
      15'b000_110100101111 : VALUE=19'b0000001_000110100000;
      15'b000_110100110000 : VALUE=19'b0000001_000110100000;
      15'b000_110100110001 : VALUE=19'b0000001_000110011111;
      15'b000_110100110010 : VALUE=19'b0000001_000110011110;
      15'b000_110100110011 : VALUE=19'b0000001_000110011110;
      15'b000_110100110100 : VALUE=19'b0000001_000110011101;
      15'b000_110100110101 : VALUE=19'b0000001_000110011100;
      15'b000_110100110110 : VALUE=19'b0000001_000110011100;
      15'b000_110100110111 : VALUE=19'b0000001_000110011011;
      15'b000_110100111000 : VALUE=19'b0000001_000110011010;
      15'b000_110100111001 : VALUE=19'b0000001_000110011010;
      15'b000_110100111010 : VALUE=19'b0000001_000110011001;
      15'b000_110100111011 : VALUE=19'b0000001_000110011000;
      15'b000_110100111100 : VALUE=19'b0000001_000110011000;
      15'b000_110100111101 : VALUE=19'b0000001_000110010111;
      15'b000_110100111110 : VALUE=19'b0000001_000110010110;
      15'b000_110100111111 : VALUE=19'b0000001_000110010110;
      15'b000_110101000000 : VALUE=19'b0000001_000110010101;
      15'b000_110101000001 : VALUE=19'b0000001_000110010100;
      15'b000_110101000010 : VALUE=19'b0000001_000110010100;
      15'b000_110101000011 : VALUE=19'b0000001_000110010011;
      15'b000_110101000100 : VALUE=19'b0000001_000110010010;
      15'b000_110101000101 : VALUE=19'b0000001_000110010010;
      15'b000_110101000110 : VALUE=19'b0000001_000110010001;
      15'b000_110101000111 : VALUE=19'b0000001_000110010000;
      15'b000_110101001000 : VALUE=19'b0000001_000110010000;
      15'b000_110101001001 : VALUE=19'b0000001_000110001111;
      15'b000_110101001010 : VALUE=19'b0000001_000110001110;
      15'b000_110101001011 : VALUE=19'b0000001_000110001110;
      15'b000_110101001100 : VALUE=19'b0000001_000110001101;
      15'b000_110101001101 : VALUE=19'b0000001_000110001100;
      15'b000_110101001110 : VALUE=19'b0000001_000110001100;
      15'b000_110101001111 : VALUE=19'b0000001_000110001011;
      15'b000_110101010000 : VALUE=19'b0000001_000110001010;
      15'b000_110101010001 : VALUE=19'b0000001_000110001010;
      15'b000_110101010010 : VALUE=19'b0000001_000110001001;
      15'b000_110101010011 : VALUE=19'b0000001_000110001000;
      15'b000_110101010100 : VALUE=19'b0000001_000110001000;
      15'b000_110101010101 : VALUE=19'b0000001_000110000111;
      15'b000_110101010110 : VALUE=19'b0000001_000110000111;
      15'b000_110101010111 : VALUE=19'b0000001_000110000110;
      15'b000_110101011000 : VALUE=19'b0000001_000110000101;
      15'b000_110101011001 : VALUE=19'b0000001_000110000101;
      15'b000_110101011010 : VALUE=19'b0000001_000110000100;
      15'b000_110101011011 : VALUE=19'b0000001_000110000011;
      15'b000_110101011100 : VALUE=19'b0000001_000110000011;
      15'b000_110101011101 : VALUE=19'b0000001_000110000010;
      15'b000_110101011110 : VALUE=19'b0000001_000110000001;
      15'b000_110101011111 : VALUE=19'b0000001_000110000001;
      15'b000_110101100000 : VALUE=19'b0000001_000110000000;
      15'b000_110101100001 : VALUE=19'b0000001_000101111111;
      15'b000_110101100010 : VALUE=19'b0000001_000101111111;
      15'b000_110101100011 : VALUE=19'b0000001_000101111110;
      15'b000_110101100100 : VALUE=19'b0000001_000101111101;
      15'b000_110101100101 : VALUE=19'b0000001_000101111101;
      15'b000_110101100110 : VALUE=19'b0000001_000101111100;
      15'b000_110101100111 : VALUE=19'b0000001_000101111011;
      15'b000_110101101000 : VALUE=19'b0000001_000101111011;
      15'b000_110101101001 : VALUE=19'b0000001_000101111010;
      15'b000_110101101010 : VALUE=19'b0000001_000101111001;
      15'b000_110101101011 : VALUE=19'b0000001_000101111001;
      15'b000_110101101100 : VALUE=19'b0000001_000101111000;
      15'b000_110101101101 : VALUE=19'b0000001_000101110111;
      15'b000_110101101110 : VALUE=19'b0000001_000101110111;
      15'b000_110101101111 : VALUE=19'b0000001_000101110110;
      15'b000_110101110000 : VALUE=19'b0000001_000101110110;
      15'b000_110101110001 : VALUE=19'b0000001_000101110101;
      15'b000_110101110010 : VALUE=19'b0000001_000101110100;
      15'b000_110101110011 : VALUE=19'b0000001_000101110100;
      15'b000_110101110100 : VALUE=19'b0000001_000101110011;
      15'b000_110101110101 : VALUE=19'b0000001_000101110010;
      15'b000_110101110110 : VALUE=19'b0000001_000101110010;
      15'b000_110101110111 : VALUE=19'b0000001_000101110001;
      15'b000_110101111000 : VALUE=19'b0000001_000101110000;
      15'b000_110101111001 : VALUE=19'b0000001_000101110000;
      15'b000_110101111010 : VALUE=19'b0000001_000101101111;
      15'b000_110101111011 : VALUE=19'b0000001_000101101110;
      15'b000_110101111100 : VALUE=19'b0000001_000101101110;
      15'b000_110101111101 : VALUE=19'b0000001_000101101101;
      15'b000_110101111110 : VALUE=19'b0000001_000101101100;
      15'b000_110101111111 : VALUE=19'b0000001_000101101100;
      15'b000_110110000000 : VALUE=19'b0000001_000101101011;
      15'b000_110110000001 : VALUE=19'b0000001_000101101011;
      15'b000_110110000010 : VALUE=19'b0000001_000101101010;
      15'b000_110110000011 : VALUE=19'b0000001_000101101001;
      15'b000_110110000100 : VALUE=19'b0000001_000101101001;
      15'b000_110110000101 : VALUE=19'b0000001_000101101000;
      15'b000_110110000110 : VALUE=19'b0000001_000101100111;
      15'b000_110110000111 : VALUE=19'b0000001_000101100111;
      15'b000_110110001000 : VALUE=19'b0000001_000101100110;
      15'b000_110110001001 : VALUE=19'b0000001_000101100101;
      15'b000_110110001010 : VALUE=19'b0000001_000101100101;
      15'b000_110110001011 : VALUE=19'b0000001_000101100100;
      15'b000_110110001100 : VALUE=19'b0000001_000101100011;
      15'b000_110110001101 : VALUE=19'b0000001_000101100011;
      15'b000_110110001110 : VALUE=19'b0000001_000101100010;
      15'b000_110110001111 : VALUE=19'b0000001_000101100010;
      15'b000_110110010000 : VALUE=19'b0000001_000101100001;
      15'b000_110110010001 : VALUE=19'b0000001_000101100000;
      15'b000_110110010010 : VALUE=19'b0000001_000101100000;
      15'b000_110110010011 : VALUE=19'b0000001_000101011111;
      15'b000_110110010100 : VALUE=19'b0000001_000101011110;
      15'b000_110110010101 : VALUE=19'b0000001_000101011110;
      15'b000_110110010110 : VALUE=19'b0000001_000101011101;
      15'b000_110110010111 : VALUE=19'b0000001_000101011100;
      15'b000_110110011000 : VALUE=19'b0000001_000101011100;
      15'b000_110110011001 : VALUE=19'b0000001_000101011011;
      15'b000_110110011010 : VALUE=19'b0000001_000101011010;
      15'b000_110110011011 : VALUE=19'b0000001_000101011010;
      15'b000_110110011100 : VALUE=19'b0000001_000101011001;
      15'b000_110110011101 : VALUE=19'b0000001_000101011001;
      15'b000_110110011110 : VALUE=19'b0000001_000101011000;
      15'b000_110110011111 : VALUE=19'b0000001_000101010111;
      15'b000_110110100000 : VALUE=19'b0000001_000101010111;
      15'b000_110110100001 : VALUE=19'b0000001_000101010110;
      15'b000_110110100010 : VALUE=19'b0000001_000101010101;
      15'b000_110110100011 : VALUE=19'b0000001_000101010101;
      15'b000_110110100100 : VALUE=19'b0000001_000101010100;
      15'b000_110110100101 : VALUE=19'b0000001_000101010011;
      15'b000_110110100110 : VALUE=19'b0000001_000101010011;
      15'b000_110110100111 : VALUE=19'b0000001_000101010010;
      15'b000_110110101000 : VALUE=19'b0000001_000101010010;
      15'b000_110110101001 : VALUE=19'b0000001_000101010001;
      15'b000_110110101010 : VALUE=19'b0000001_000101010000;
      15'b000_110110101011 : VALUE=19'b0000001_000101010000;
      15'b000_110110101100 : VALUE=19'b0000001_000101001111;
      15'b000_110110101101 : VALUE=19'b0000001_000101001110;
      15'b000_110110101110 : VALUE=19'b0000001_000101001110;
      15'b000_110110101111 : VALUE=19'b0000001_000101001101;
      15'b000_110110110000 : VALUE=19'b0000001_000101001101;
      15'b000_110110110001 : VALUE=19'b0000001_000101001100;
      15'b000_110110110010 : VALUE=19'b0000001_000101001011;
      15'b000_110110110011 : VALUE=19'b0000001_000101001011;
      15'b000_110110110100 : VALUE=19'b0000001_000101001010;
      15'b000_110110110101 : VALUE=19'b0000001_000101001001;
      15'b000_110110110110 : VALUE=19'b0000001_000101001001;
      15'b000_110110110111 : VALUE=19'b0000001_000101001000;
      15'b000_110110111000 : VALUE=19'b0000001_000101000111;
      15'b000_110110111001 : VALUE=19'b0000001_000101000111;
      15'b000_110110111010 : VALUE=19'b0000001_000101000110;
      15'b000_110110111011 : VALUE=19'b0000001_000101000110;
      15'b000_110110111100 : VALUE=19'b0000001_000101000101;
      15'b000_110110111101 : VALUE=19'b0000001_000101000100;
      15'b000_110110111110 : VALUE=19'b0000001_000101000100;
      15'b000_110110111111 : VALUE=19'b0000001_000101000011;
      15'b000_110111000000 : VALUE=19'b0000001_000101000010;
      15'b000_110111000001 : VALUE=19'b0000001_000101000010;
      15'b000_110111000010 : VALUE=19'b0000001_000101000001;
      15'b000_110111000011 : VALUE=19'b0000001_000101000001;
      15'b000_110111000100 : VALUE=19'b0000001_000101000000;
      15'b000_110111000101 : VALUE=19'b0000001_000100111111;
      15'b000_110111000110 : VALUE=19'b0000001_000100111111;
      15'b000_110111000111 : VALUE=19'b0000001_000100111110;
      15'b000_110111001000 : VALUE=19'b0000001_000100111101;
      15'b000_110111001001 : VALUE=19'b0000001_000100111101;
      15'b000_110111001010 : VALUE=19'b0000001_000100111100;
      15'b000_110111001011 : VALUE=19'b0000001_000100111100;
      15'b000_110111001100 : VALUE=19'b0000001_000100111011;
      15'b000_110111001101 : VALUE=19'b0000001_000100111010;
      15'b000_110111001110 : VALUE=19'b0000001_000100111010;
      15'b000_110111001111 : VALUE=19'b0000001_000100111001;
      15'b000_110111010000 : VALUE=19'b0000001_000100111000;
      15'b000_110111010001 : VALUE=19'b0000001_000100111000;
      15'b000_110111010010 : VALUE=19'b0000001_000100110111;
      15'b000_110111010011 : VALUE=19'b0000001_000100110111;
      15'b000_110111010100 : VALUE=19'b0000001_000100110110;
      15'b000_110111010101 : VALUE=19'b0000001_000100110101;
      15'b000_110111010110 : VALUE=19'b0000001_000100110101;
      15'b000_110111010111 : VALUE=19'b0000001_000100110100;
      15'b000_110111011000 : VALUE=19'b0000001_000100110011;
      15'b000_110111011001 : VALUE=19'b0000001_000100110011;
      15'b000_110111011010 : VALUE=19'b0000001_000100110010;
      15'b000_110111011011 : VALUE=19'b0000001_000100110010;
      15'b000_110111011100 : VALUE=19'b0000001_000100110001;
      15'b000_110111011101 : VALUE=19'b0000001_000100110000;
      15'b000_110111011110 : VALUE=19'b0000001_000100110000;
      15'b000_110111011111 : VALUE=19'b0000001_000100101111;
      15'b000_110111100000 : VALUE=19'b0000001_000100101110;
      15'b000_110111100001 : VALUE=19'b0000001_000100101110;
      15'b000_110111100010 : VALUE=19'b0000001_000100101101;
      15'b000_110111100011 : VALUE=19'b0000001_000100101101;
      15'b000_110111100100 : VALUE=19'b0000001_000100101100;
      15'b000_110111100101 : VALUE=19'b0000001_000100101011;
      15'b000_110111100110 : VALUE=19'b0000001_000100101011;
      15'b000_110111100111 : VALUE=19'b0000001_000100101010;
      15'b000_110111101000 : VALUE=19'b0000001_000100101010;
      15'b000_110111101001 : VALUE=19'b0000001_000100101001;
      15'b000_110111101010 : VALUE=19'b0000001_000100101000;
      15'b000_110111101011 : VALUE=19'b0000001_000100101000;
      15'b000_110111101100 : VALUE=19'b0000001_000100100111;
      15'b000_110111101101 : VALUE=19'b0000001_000100100110;
      15'b000_110111101110 : VALUE=19'b0000001_000100100110;
      15'b000_110111101111 : VALUE=19'b0000001_000100100101;
      15'b000_110111110000 : VALUE=19'b0000001_000100100101;
      15'b000_110111110001 : VALUE=19'b0000001_000100100100;
      15'b000_110111110010 : VALUE=19'b0000001_000100100011;
      15'b000_110111110011 : VALUE=19'b0000001_000100100011;
      15'b000_110111110100 : VALUE=19'b0000001_000100100010;
      15'b000_110111110101 : VALUE=19'b0000001_000100100010;
      15'b000_110111110110 : VALUE=19'b0000001_000100100001;
      15'b000_110111110111 : VALUE=19'b0000001_000100100000;
      15'b000_110111111000 : VALUE=19'b0000001_000100100000;
      15'b000_110111111001 : VALUE=19'b0000001_000100011111;
      15'b000_110111111010 : VALUE=19'b0000001_000100011110;
      15'b000_110111111011 : VALUE=19'b0000001_000100011110;
      15'b000_110111111100 : VALUE=19'b0000001_000100011101;
      15'b000_110111111101 : VALUE=19'b0000001_000100011101;
      15'b000_110111111110 : VALUE=19'b0000001_000100011100;
      15'b000_110111111111 : VALUE=19'b0000001_000100011011;
      15'b000_111000000000 : VALUE=19'b0000001_000100011011;
      15'b000_111000000001 : VALUE=19'b0000001_000100011010;
      15'b000_111000000010 : VALUE=19'b0000001_000100011010;
      15'b000_111000000011 : VALUE=19'b0000001_000100011001;
      15'b000_111000000100 : VALUE=19'b0000001_000100011000;
      15'b000_111000000101 : VALUE=19'b0000001_000100011000;
      15'b000_111000000110 : VALUE=19'b0000001_000100010111;
      15'b000_111000000111 : VALUE=19'b0000001_000100010111;
      15'b000_111000001000 : VALUE=19'b0000001_000100010110;
      15'b000_111000001001 : VALUE=19'b0000001_000100010101;
      15'b000_111000001010 : VALUE=19'b0000001_000100010101;
      15'b000_111000001011 : VALUE=19'b0000001_000100010100;
      15'b000_111000001100 : VALUE=19'b0000001_000100010011;
      15'b000_111000001101 : VALUE=19'b0000001_000100010011;
      15'b000_111000001110 : VALUE=19'b0000001_000100010010;
      15'b000_111000001111 : VALUE=19'b0000001_000100010010;
      15'b000_111000010000 : VALUE=19'b0000001_000100010001;
      15'b000_111000010001 : VALUE=19'b0000001_000100010000;
      15'b000_111000010010 : VALUE=19'b0000001_000100010000;
      15'b000_111000010011 : VALUE=19'b0000001_000100001111;
      15'b000_111000010100 : VALUE=19'b0000001_000100001111;
      15'b000_111000010101 : VALUE=19'b0000001_000100001110;
      15'b000_111000010110 : VALUE=19'b0000001_000100001101;
      15'b000_111000010111 : VALUE=19'b0000001_000100001101;
      15'b000_111000011000 : VALUE=19'b0000001_000100001100;
      15'b000_111000011001 : VALUE=19'b0000001_000100001100;
      15'b000_111000011010 : VALUE=19'b0000001_000100001011;
      15'b000_111000011011 : VALUE=19'b0000001_000100001010;
      15'b000_111000011100 : VALUE=19'b0000001_000100001010;
      15'b000_111000011101 : VALUE=19'b0000001_000100001001;
      15'b000_111000011110 : VALUE=19'b0000001_000100001001;
      15'b000_111000011111 : VALUE=19'b0000001_000100001000;
      15'b000_111000100000 : VALUE=19'b0000001_000100000111;
      15'b000_111000100001 : VALUE=19'b0000001_000100000111;
      15'b000_111000100010 : VALUE=19'b0000001_000100000110;
      15'b000_111000100011 : VALUE=19'b0000001_000100000110;
      15'b000_111000100100 : VALUE=19'b0000001_000100000101;
      15'b000_111000100101 : VALUE=19'b0000001_000100000100;
      15'b000_111000100110 : VALUE=19'b0000001_000100000100;
      15'b000_111000100111 : VALUE=19'b0000001_000100000011;
      15'b000_111000101000 : VALUE=19'b0000001_000100000011;
      15'b000_111000101001 : VALUE=19'b0000001_000100000010;
      15'b000_111000101010 : VALUE=19'b0000001_000100000001;
      15'b000_111000101011 : VALUE=19'b0000001_000100000001;
      15'b000_111000101100 : VALUE=19'b0000001_000100000000;
      15'b000_111000101101 : VALUE=19'b0000001_000100000000;
      15'b000_111000101110 : VALUE=19'b0000001_000011111111;
      15'b000_111000101111 : VALUE=19'b0000001_000011111110;
      15'b000_111000110000 : VALUE=19'b0000001_000011111110;
      15'b000_111000110001 : VALUE=19'b0000001_000011111101;
      15'b000_111000110010 : VALUE=19'b0000001_000011111101;
      15'b000_111000110011 : VALUE=19'b0000001_000011111100;
      15'b000_111000110100 : VALUE=19'b0000001_000011111011;
      15'b000_111000110101 : VALUE=19'b0000001_000011111011;
      15'b000_111000110110 : VALUE=19'b0000001_000011111010;
      15'b000_111000110111 : VALUE=19'b0000001_000011111010;
      15'b000_111000111000 : VALUE=19'b0000001_000011111001;
      15'b000_111000111001 : VALUE=19'b0000001_000011111000;
      15'b000_111000111010 : VALUE=19'b0000001_000011111000;
      15'b000_111000111011 : VALUE=19'b0000001_000011110111;
      15'b000_111000111100 : VALUE=19'b0000001_000011110111;
      15'b000_111000111101 : VALUE=19'b0000001_000011110110;
      15'b000_111000111110 : VALUE=19'b0000001_000011110101;
      15'b000_111000111111 : VALUE=19'b0000001_000011110101;
      15'b000_111001000000 : VALUE=19'b0000001_000011110100;
      15'b000_111001000001 : VALUE=19'b0000001_000011110100;
      15'b000_111001000010 : VALUE=19'b0000001_000011110011;
      15'b000_111001000011 : VALUE=19'b0000001_000011110010;
      15'b000_111001000100 : VALUE=19'b0000001_000011110010;
      15'b000_111001000101 : VALUE=19'b0000001_000011110001;
      15'b000_111001000110 : VALUE=19'b0000001_000011110001;
      15'b000_111001000111 : VALUE=19'b0000001_000011110000;
      15'b000_111001001000 : VALUE=19'b0000001_000011101111;
      15'b000_111001001001 : VALUE=19'b0000001_000011101111;
      15'b000_111001001010 : VALUE=19'b0000001_000011101110;
      15'b000_111001001011 : VALUE=19'b0000001_000011101110;
      15'b000_111001001100 : VALUE=19'b0000001_000011101101;
      15'b000_111001001101 : VALUE=19'b0000001_000011101101;
      15'b000_111001001110 : VALUE=19'b0000001_000011101100;
      15'b000_111001001111 : VALUE=19'b0000001_000011101011;
      15'b000_111001010000 : VALUE=19'b0000001_000011101011;
      15'b000_111001010001 : VALUE=19'b0000001_000011101010;
      15'b000_111001010010 : VALUE=19'b0000001_000011101010;
      15'b000_111001010011 : VALUE=19'b0000001_000011101001;
      15'b000_111001010100 : VALUE=19'b0000001_000011101000;
      15'b000_111001010101 : VALUE=19'b0000001_000011101000;
      15'b000_111001010110 : VALUE=19'b0000001_000011100111;
      15'b000_111001010111 : VALUE=19'b0000001_000011100111;
      15'b000_111001011000 : VALUE=19'b0000001_000011100110;
      15'b000_111001011001 : VALUE=19'b0000001_000011100101;
      15'b000_111001011010 : VALUE=19'b0000001_000011100101;
      15'b000_111001011011 : VALUE=19'b0000001_000011100100;
      15'b000_111001011100 : VALUE=19'b0000001_000011100100;
      15'b000_111001011101 : VALUE=19'b0000001_000011100011;
      15'b000_111001011110 : VALUE=19'b0000001_000011100010;
      15'b000_111001011111 : VALUE=19'b0000001_000011100010;
      15'b000_111001100000 : VALUE=19'b0000001_000011100001;
      15'b000_111001100001 : VALUE=19'b0000001_000011100001;
      15'b000_111001100010 : VALUE=19'b0000001_000011100000;
      15'b000_111001100011 : VALUE=19'b0000001_000011100000;
      15'b000_111001100100 : VALUE=19'b0000001_000011011111;
      15'b000_111001100101 : VALUE=19'b0000001_000011011110;
      15'b000_111001100110 : VALUE=19'b0000001_000011011110;
      15'b000_111001100111 : VALUE=19'b0000001_000011011101;
      15'b000_111001101000 : VALUE=19'b0000001_000011011101;
      15'b000_111001101001 : VALUE=19'b0000001_000011011100;
      15'b000_111001101010 : VALUE=19'b0000001_000011011011;
      15'b000_111001101011 : VALUE=19'b0000001_000011011011;
      15'b000_111001101100 : VALUE=19'b0000001_000011011010;
      15'b000_111001101101 : VALUE=19'b0000001_000011011010;
      15'b000_111001101110 : VALUE=19'b0000001_000011011001;
      15'b000_111001101111 : VALUE=19'b0000001_000011011001;
      15'b000_111001110000 : VALUE=19'b0000001_000011011000;
      15'b000_111001110001 : VALUE=19'b0000001_000011010111;
      15'b000_111001110010 : VALUE=19'b0000001_000011010111;
      15'b000_111001110011 : VALUE=19'b0000001_000011010110;
      15'b000_111001110100 : VALUE=19'b0000001_000011010110;
      15'b000_111001110101 : VALUE=19'b0000001_000011010101;
      15'b000_111001110110 : VALUE=19'b0000001_000011010100;
      15'b000_111001110111 : VALUE=19'b0000001_000011010100;
      15'b000_111001111000 : VALUE=19'b0000001_000011010011;
      15'b000_111001111001 : VALUE=19'b0000001_000011010011;
      15'b000_111001111010 : VALUE=19'b0000001_000011010010;
      15'b000_111001111011 : VALUE=19'b0000001_000011010010;
      15'b000_111001111100 : VALUE=19'b0000001_000011010001;
      15'b000_111001111101 : VALUE=19'b0000001_000011010000;
      15'b000_111001111110 : VALUE=19'b0000001_000011010000;
      15'b000_111001111111 : VALUE=19'b0000001_000011001111;
      15'b000_111010000000 : VALUE=19'b0000001_000011001111;
      15'b000_111010000001 : VALUE=19'b0000001_000011001110;
      15'b000_111010000010 : VALUE=19'b0000001_000011001101;
      15'b000_111010000011 : VALUE=19'b0000001_000011001101;
      15'b000_111010000100 : VALUE=19'b0000001_000011001100;
      15'b000_111010000101 : VALUE=19'b0000001_000011001100;
      15'b000_111010000110 : VALUE=19'b0000001_000011001011;
      15'b000_111010000111 : VALUE=19'b0000001_000011001011;
      15'b000_111010001000 : VALUE=19'b0000001_000011001010;
      15'b000_111010001001 : VALUE=19'b0000001_000011001001;
      15'b000_111010001010 : VALUE=19'b0000001_000011001001;
      15'b000_111010001011 : VALUE=19'b0000001_000011001000;
      15'b000_111010001100 : VALUE=19'b0000001_000011001000;
      15'b000_111010001101 : VALUE=19'b0000001_000011000111;
      15'b000_111010001110 : VALUE=19'b0000001_000011000111;
      15'b000_111010001111 : VALUE=19'b0000001_000011000110;
      15'b000_111010010000 : VALUE=19'b0000001_000011000101;
      15'b000_111010010001 : VALUE=19'b0000001_000011000101;
      15'b000_111010010010 : VALUE=19'b0000001_000011000100;
      15'b000_111010010011 : VALUE=19'b0000001_000011000100;
      15'b000_111010010100 : VALUE=19'b0000001_000011000011;
      15'b000_111010010101 : VALUE=19'b0000001_000011000011;
      15'b000_111010010110 : VALUE=19'b0000001_000011000010;
      15'b000_111010010111 : VALUE=19'b0000001_000011000001;
      15'b000_111010011000 : VALUE=19'b0000001_000011000001;
      15'b000_111010011001 : VALUE=19'b0000001_000011000000;
      15'b000_111010011010 : VALUE=19'b0000001_000011000000;
      15'b000_111010011011 : VALUE=19'b0000001_000010111111;
      15'b000_111010011100 : VALUE=19'b0000001_000010111111;
      15'b000_111010011101 : VALUE=19'b0000001_000010111110;
      15'b000_111010011110 : VALUE=19'b0000001_000010111101;
      15'b000_111010011111 : VALUE=19'b0000001_000010111101;
      15'b000_111010100000 : VALUE=19'b0000001_000010111100;
      15'b000_111010100001 : VALUE=19'b0000001_000010111100;
      15'b000_111010100010 : VALUE=19'b0000001_000010111011;
      15'b000_111010100011 : VALUE=19'b0000001_000010111011;
      15'b000_111010100100 : VALUE=19'b0000001_000010111010;
      15'b000_111010100101 : VALUE=19'b0000001_000010111001;
      15'b000_111010100110 : VALUE=19'b0000001_000010111001;
      15'b000_111010100111 : VALUE=19'b0000001_000010111000;
      15'b000_111010101000 : VALUE=19'b0000001_000010111000;
      15'b000_111010101001 : VALUE=19'b0000001_000010110111;
      15'b000_111010101010 : VALUE=19'b0000001_000010110111;
      15'b000_111010101011 : VALUE=19'b0000001_000010110110;
      15'b000_111010101100 : VALUE=19'b0000001_000010110101;
      15'b000_111010101101 : VALUE=19'b0000001_000010110101;
      15'b000_111010101110 : VALUE=19'b0000001_000010110100;
      15'b000_111010101111 : VALUE=19'b0000001_000010110100;
      15'b000_111010110000 : VALUE=19'b0000001_000010110011;
      15'b000_111010110001 : VALUE=19'b0000001_000010110011;
      15'b000_111010110010 : VALUE=19'b0000001_000010110010;
      15'b000_111010110011 : VALUE=19'b0000001_000010110001;
      15'b000_111010110100 : VALUE=19'b0000001_000010110001;
      15'b000_111010110101 : VALUE=19'b0000001_000010110000;
      15'b000_111010110110 : VALUE=19'b0000001_000010110000;
      15'b000_111010110111 : VALUE=19'b0000001_000010101111;
      15'b000_111010111000 : VALUE=19'b0000001_000010101111;
      15'b000_111010111001 : VALUE=19'b0000001_000010101110;
      15'b000_111010111010 : VALUE=19'b0000001_000010101101;
      15'b000_111010111011 : VALUE=19'b0000001_000010101101;
      15'b000_111010111100 : VALUE=19'b0000001_000010101100;
      15'b000_111010111101 : VALUE=19'b0000001_000010101100;
      15'b000_111010111110 : VALUE=19'b0000001_000010101011;
      15'b000_111010111111 : VALUE=19'b0000001_000010101011;
      15'b000_111011000000 : VALUE=19'b0000001_000010101010;
      15'b000_111011000001 : VALUE=19'b0000001_000010101001;
      15'b000_111011000010 : VALUE=19'b0000001_000010101001;
      15'b000_111011000011 : VALUE=19'b0000001_000010101000;
      15'b000_111011000100 : VALUE=19'b0000001_000010101000;
      15'b000_111011000101 : VALUE=19'b0000001_000010100111;
      15'b000_111011000110 : VALUE=19'b0000001_000010100111;
      15'b000_111011000111 : VALUE=19'b0000001_000010100110;
      15'b000_111011001000 : VALUE=19'b0000001_000010100110;
      15'b000_111011001001 : VALUE=19'b0000001_000010100101;
      15'b000_111011001010 : VALUE=19'b0000001_000010100100;
      15'b000_111011001011 : VALUE=19'b0000001_000010100100;
      15'b000_111011001100 : VALUE=19'b0000001_000010100011;
      15'b000_111011001101 : VALUE=19'b0000001_000010100011;
      15'b000_111011001110 : VALUE=19'b0000001_000010100010;
      15'b000_111011001111 : VALUE=19'b0000001_000010100010;
      15'b000_111011010000 : VALUE=19'b0000001_000010100001;
      15'b000_111011010001 : VALUE=19'b0000001_000010100000;
      15'b000_111011010010 : VALUE=19'b0000001_000010100000;
      15'b000_111011010011 : VALUE=19'b0000001_000010011111;
      15'b000_111011010100 : VALUE=19'b0000001_000010011111;
      15'b000_111011010101 : VALUE=19'b0000001_000010011110;
      15'b000_111011010110 : VALUE=19'b0000001_000010011110;
      15'b000_111011010111 : VALUE=19'b0000001_000010011101;
      15'b000_111011011000 : VALUE=19'b0000001_000010011101;
      15'b000_111011011001 : VALUE=19'b0000001_000010011100;
      15'b000_111011011010 : VALUE=19'b0000001_000010011011;
      15'b000_111011011011 : VALUE=19'b0000001_000010011011;
      15'b000_111011011100 : VALUE=19'b0000001_000010011010;
      15'b000_111011011101 : VALUE=19'b0000001_000010011010;
      15'b000_111011011110 : VALUE=19'b0000001_000010011001;
      15'b000_111011011111 : VALUE=19'b0000001_000010011001;
      15'b000_111011100000 : VALUE=19'b0000001_000010011000;
      15'b000_111011100001 : VALUE=19'b0000001_000010011000;
      15'b000_111011100010 : VALUE=19'b0000001_000010010111;
      15'b000_111011100011 : VALUE=19'b0000001_000010010110;
      15'b000_111011100100 : VALUE=19'b0000001_000010010110;
      15'b000_111011100101 : VALUE=19'b0000001_000010010101;
      15'b000_111011100110 : VALUE=19'b0000001_000010010101;
      15'b000_111011100111 : VALUE=19'b0000001_000010010100;
      15'b000_111011101000 : VALUE=19'b0000001_000010010100;
      15'b000_111011101001 : VALUE=19'b0000001_000010010011;
      15'b000_111011101010 : VALUE=19'b0000001_000010010011;
      15'b000_111011101011 : VALUE=19'b0000001_000010010010;
      15'b000_111011101100 : VALUE=19'b0000001_000010010001;
      15'b000_111011101101 : VALUE=19'b0000001_000010010001;
      15'b000_111011101110 : VALUE=19'b0000001_000010010000;
      15'b000_111011101111 : VALUE=19'b0000001_000010010000;
      15'b000_111011110000 : VALUE=19'b0000001_000010001111;
      15'b000_111011110001 : VALUE=19'b0000001_000010001111;
      15'b000_111011110010 : VALUE=19'b0000001_000010001110;
      15'b000_111011110011 : VALUE=19'b0000001_000010001110;
      15'b000_111011110100 : VALUE=19'b0000001_000010001101;
      15'b000_111011110101 : VALUE=19'b0000001_000010001100;
      15'b000_111011110110 : VALUE=19'b0000001_000010001100;
      15'b000_111011110111 : VALUE=19'b0000001_000010001011;
      15'b000_111011111000 : VALUE=19'b0000001_000010001011;
      15'b000_111011111001 : VALUE=19'b0000001_000010001010;
      15'b000_111011111010 : VALUE=19'b0000001_000010001010;
      15'b000_111011111011 : VALUE=19'b0000001_000010001001;
      15'b000_111011111100 : VALUE=19'b0000001_000010001001;
      15'b000_111011111101 : VALUE=19'b0000001_000010001000;
      15'b000_111011111110 : VALUE=19'b0000001_000010000111;
      15'b000_111011111111 : VALUE=19'b0000001_000010000111;
      15'b000_111100000000 : VALUE=19'b0000001_000010000110;
      15'b000_111100000001 : VALUE=19'b0000001_000010000110;
      15'b000_111100000010 : VALUE=19'b0000001_000010000101;
      15'b000_111100000011 : VALUE=19'b0000001_000010000101;
      15'b000_111100000100 : VALUE=19'b0000001_000010000100;
      15'b000_111100000101 : VALUE=19'b0000001_000010000100;
      15'b000_111100000110 : VALUE=19'b0000001_000010000011;
      15'b000_111100000111 : VALUE=19'b0000001_000010000010;
      15'b000_111100001000 : VALUE=19'b0000001_000010000010;
      15'b000_111100001001 : VALUE=19'b0000001_000010000001;
      15'b000_111100001010 : VALUE=19'b0000001_000010000001;
      15'b000_111100001011 : VALUE=19'b0000001_000010000000;
      15'b000_111100001100 : VALUE=19'b0000001_000010000000;
      15'b000_111100001101 : VALUE=19'b0000001_000001111111;
      15'b000_111100001110 : VALUE=19'b0000001_000001111111;
      15'b000_111100001111 : VALUE=19'b0000001_000001111110;
      15'b000_111100010000 : VALUE=19'b0000001_000001111110;
      15'b000_111100010001 : VALUE=19'b0000001_000001111101;
      15'b000_111100010010 : VALUE=19'b0000001_000001111100;
      15'b000_111100010011 : VALUE=19'b0000001_000001111100;
      15'b000_111100010100 : VALUE=19'b0000001_000001111011;
      15'b000_111100010101 : VALUE=19'b0000001_000001111011;
      15'b000_111100010110 : VALUE=19'b0000001_000001111010;
      15'b000_111100010111 : VALUE=19'b0000001_000001111010;
      15'b000_111100011000 : VALUE=19'b0000001_000001111001;
      15'b000_111100011001 : VALUE=19'b0000001_000001111001;
      15'b000_111100011010 : VALUE=19'b0000001_000001111000;
      15'b000_111100011011 : VALUE=19'b0000001_000001111000;
      15'b000_111100011100 : VALUE=19'b0000001_000001110111;
      15'b000_111100011101 : VALUE=19'b0000001_000001110110;
      15'b000_111100011110 : VALUE=19'b0000001_000001110110;
      15'b000_111100011111 : VALUE=19'b0000001_000001110101;
      15'b000_111100100000 : VALUE=19'b0000001_000001110101;
      15'b000_111100100001 : VALUE=19'b0000001_000001110100;
      15'b000_111100100010 : VALUE=19'b0000001_000001110100;
      15'b000_111100100011 : VALUE=19'b0000001_000001110011;
      15'b000_111100100100 : VALUE=19'b0000001_000001110011;
      15'b000_111100100101 : VALUE=19'b0000001_000001110010;
      15'b000_111100100110 : VALUE=19'b0000001_000001110010;
      15'b000_111100100111 : VALUE=19'b0000001_000001110001;
      15'b000_111100101000 : VALUE=19'b0000001_000001110000;
      15'b000_111100101001 : VALUE=19'b0000001_000001110000;
      15'b000_111100101010 : VALUE=19'b0000001_000001101111;
      15'b000_111100101011 : VALUE=19'b0000001_000001101111;
      15'b000_111100101100 : VALUE=19'b0000001_000001101110;
      15'b000_111100101101 : VALUE=19'b0000001_000001101110;
      15'b000_111100101110 : VALUE=19'b0000001_000001101101;
      15'b000_111100101111 : VALUE=19'b0000001_000001101101;
      15'b000_111100110000 : VALUE=19'b0000001_000001101100;
      15'b000_111100110001 : VALUE=19'b0000001_000001101100;
      15'b000_111100110010 : VALUE=19'b0000001_000001101011;
      15'b000_111100110011 : VALUE=19'b0000001_000001101011;
      15'b000_111100110100 : VALUE=19'b0000001_000001101010;
      15'b000_111100110101 : VALUE=19'b0000001_000001101001;
      15'b000_111100110110 : VALUE=19'b0000001_000001101001;
      15'b000_111100110111 : VALUE=19'b0000001_000001101000;
      15'b000_111100111000 : VALUE=19'b0000001_000001101000;
      15'b000_111100111001 : VALUE=19'b0000001_000001100111;
      15'b000_111100111010 : VALUE=19'b0000001_000001100111;
      15'b000_111100111011 : VALUE=19'b0000001_000001100110;
      15'b000_111100111100 : VALUE=19'b0000001_000001100110;
      15'b000_111100111101 : VALUE=19'b0000001_000001100101;
      15'b000_111100111110 : VALUE=19'b0000001_000001100101;
      15'b000_111100111111 : VALUE=19'b0000001_000001100100;
      15'b000_111101000000 : VALUE=19'b0000001_000001100100;
      15'b000_111101000001 : VALUE=19'b0000001_000001100011;
      15'b000_111101000010 : VALUE=19'b0000001_000001100010;
      15'b000_111101000011 : VALUE=19'b0000001_000001100010;
      15'b000_111101000100 : VALUE=19'b0000001_000001100001;
      15'b000_111101000101 : VALUE=19'b0000001_000001100001;
      15'b000_111101000110 : VALUE=19'b0000001_000001100000;
      15'b000_111101000111 : VALUE=19'b0000001_000001100000;
      15'b000_111101001000 : VALUE=19'b0000001_000001011111;
      15'b000_111101001001 : VALUE=19'b0000001_000001011111;
      15'b000_111101001010 : VALUE=19'b0000001_000001011110;
      15'b000_111101001011 : VALUE=19'b0000001_000001011110;
      15'b000_111101001100 : VALUE=19'b0000001_000001011101;
      15'b000_111101001101 : VALUE=19'b0000001_000001011101;
      15'b000_111101001110 : VALUE=19'b0000001_000001011100;
      15'b000_111101001111 : VALUE=19'b0000001_000001011011;
      15'b000_111101010000 : VALUE=19'b0000001_000001011011;
      15'b000_111101010001 : VALUE=19'b0000001_000001011010;
      15'b000_111101010010 : VALUE=19'b0000001_000001011010;
      15'b000_111101010011 : VALUE=19'b0000001_000001011001;
      15'b000_111101010100 : VALUE=19'b0000001_000001011001;
      15'b000_111101010101 : VALUE=19'b0000001_000001011000;
      15'b000_111101010110 : VALUE=19'b0000001_000001011000;
      15'b000_111101010111 : VALUE=19'b0000001_000001010111;
      15'b000_111101011000 : VALUE=19'b0000001_000001010111;
      15'b000_111101011001 : VALUE=19'b0000001_000001010110;
      15'b000_111101011010 : VALUE=19'b0000001_000001010110;
      15'b000_111101011011 : VALUE=19'b0000001_000001010101;
      15'b000_111101011100 : VALUE=19'b0000001_000001010101;
      15'b000_111101011101 : VALUE=19'b0000001_000001010100;
      15'b000_111101011110 : VALUE=19'b0000001_000001010011;
      15'b000_111101011111 : VALUE=19'b0000001_000001010011;
      15'b000_111101100000 : VALUE=19'b0000001_000001010010;
      15'b000_111101100001 : VALUE=19'b0000001_000001010010;
      15'b000_111101100010 : VALUE=19'b0000001_000001010001;
      15'b000_111101100011 : VALUE=19'b0000001_000001010001;
      15'b000_111101100100 : VALUE=19'b0000001_000001010000;
      15'b000_111101100101 : VALUE=19'b0000001_000001010000;
      15'b000_111101100110 : VALUE=19'b0000001_000001001111;
      15'b000_111101100111 : VALUE=19'b0000001_000001001111;
      15'b000_111101101000 : VALUE=19'b0000001_000001001110;
      15'b000_111101101001 : VALUE=19'b0000001_000001001110;
      15'b000_111101101010 : VALUE=19'b0000001_000001001101;
      15'b000_111101101011 : VALUE=19'b0000001_000001001101;
      15'b000_111101101100 : VALUE=19'b0000001_000001001100;
      15'b000_111101101101 : VALUE=19'b0000001_000001001100;
      15'b000_111101101110 : VALUE=19'b0000001_000001001011;
      15'b000_111101101111 : VALUE=19'b0000001_000001001010;
      15'b000_111101110000 : VALUE=19'b0000001_000001001010;
      15'b000_111101110001 : VALUE=19'b0000001_000001001001;
      15'b000_111101110010 : VALUE=19'b0000001_000001001001;
      15'b000_111101110011 : VALUE=19'b0000001_000001001000;
      15'b000_111101110100 : VALUE=19'b0000001_000001001000;
      15'b000_111101110101 : VALUE=19'b0000001_000001000111;
      15'b000_111101110110 : VALUE=19'b0000001_000001000111;
      15'b000_111101110111 : VALUE=19'b0000001_000001000110;
      15'b000_111101111000 : VALUE=19'b0000001_000001000110;
      15'b000_111101111001 : VALUE=19'b0000001_000001000101;
      15'b000_111101111010 : VALUE=19'b0000001_000001000101;
      15'b000_111101111011 : VALUE=19'b0000001_000001000100;
      15'b000_111101111100 : VALUE=19'b0000001_000001000100;
      15'b000_111101111101 : VALUE=19'b0000001_000001000011;
      15'b000_111101111110 : VALUE=19'b0000001_000001000011;
      15'b000_111101111111 : VALUE=19'b0000001_000001000010;
      15'b000_111110000000 : VALUE=19'b0000001_000001000010;
      15'b000_111110000001 : VALUE=19'b0000001_000001000001;
      15'b000_111110000010 : VALUE=19'b0000001_000001000000;
      15'b000_111110000011 : VALUE=19'b0000001_000001000000;
      15'b000_111110000100 : VALUE=19'b0000001_000000111111;
      15'b000_111110000101 : VALUE=19'b0000001_000000111111;
      15'b000_111110000110 : VALUE=19'b0000001_000000111110;
      15'b000_111110000111 : VALUE=19'b0000001_000000111110;
      15'b000_111110001000 : VALUE=19'b0000001_000000111101;
      15'b000_111110001001 : VALUE=19'b0000001_000000111101;
      15'b000_111110001010 : VALUE=19'b0000001_000000111100;
      15'b000_111110001011 : VALUE=19'b0000001_000000111100;
      15'b000_111110001100 : VALUE=19'b0000001_000000111011;
      15'b000_111110001101 : VALUE=19'b0000001_000000111011;
      15'b000_111110001110 : VALUE=19'b0000001_000000111010;
      15'b000_111110001111 : VALUE=19'b0000001_000000111010;
      15'b000_111110010000 : VALUE=19'b0000001_000000111001;
      15'b000_111110010001 : VALUE=19'b0000001_000000111001;
      15'b000_111110010010 : VALUE=19'b0000001_000000111000;
      15'b000_111110010011 : VALUE=19'b0000001_000000111000;
      15'b000_111110010100 : VALUE=19'b0000001_000000110111;
      15'b000_111110010101 : VALUE=19'b0000001_000000110111;
      15'b000_111110010110 : VALUE=19'b0000001_000000110110;
      15'b000_111110010111 : VALUE=19'b0000001_000000110110;
      15'b000_111110011000 : VALUE=19'b0000001_000000110101;
      15'b000_111110011001 : VALUE=19'b0000001_000000110100;
      15'b000_111110011010 : VALUE=19'b0000001_000000110100;
      15'b000_111110011011 : VALUE=19'b0000001_000000110011;
      15'b000_111110011100 : VALUE=19'b0000001_000000110011;
      15'b000_111110011101 : VALUE=19'b0000001_000000110010;
      15'b000_111110011110 : VALUE=19'b0000001_000000110010;
      15'b000_111110011111 : VALUE=19'b0000001_000000110001;
      15'b000_111110100000 : VALUE=19'b0000001_000000110001;
      15'b000_111110100001 : VALUE=19'b0000001_000000110000;
      15'b000_111110100010 : VALUE=19'b0000001_000000110000;
      15'b000_111110100011 : VALUE=19'b0000001_000000101111;
      15'b000_111110100100 : VALUE=19'b0000001_000000101111;
      15'b000_111110100101 : VALUE=19'b0000001_000000101110;
      15'b000_111110100110 : VALUE=19'b0000001_000000101110;
      15'b000_111110100111 : VALUE=19'b0000001_000000101101;
      15'b000_111110101000 : VALUE=19'b0000001_000000101101;
      15'b000_111110101001 : VALUE=19'b0000001_000000101100;
      15'b000_111110101010 : VALUE=19'b0000001_000000101100;
      15'b000_111110101011 : VALUE=19'b0000001_000000101011;
      15'b000_111110101100 : VALUE=19'b0000001_000000101011;
      15'b000_111110101101 : VALUE=19'b0000001_000000101010;
      15'b000_111110101110 : VALUE=19'b0000001_000000101010;
      15'b000_111110101111 : VALUE=19'b0000001_000000101001;
      15'b000_111110110000 : VALUE=19'b0000001_000000101001;
      15'b000_111110110001 : VALUE=19'b0000001_000000101000;
      15'b000_111110110010 : VALUE=19'b0000001_000000101000;
      15'b000_111110110011 : VALUE=19'b0000001_000000100111;
      15'b000_111110110100 : VALUE=19'b0000001_000000100111;
      15'b000_111110110101 : VALUE=19'b0000001_000000100110;
      15'b000_111110110110 : VALUE=19'b0000001_000000100110;
      15'b000_111110110111 : VALUE=19'b0000001_000000100101;
      15'b000_111110111000 : VALUE=19'b0000001_000000100100;
      15'b000_111110111001 : VALUE=19'b0000001_000000100100;
      15'b000_111110111010 : VALUE=19'b0000001_000000100011;
      15'b000_111110111011 : VALUE=19'b0000001_000000100011;
      15'b000_111110111100 : VALUE=19'b0000001_000000100010;
      15'b000_111110111101 : VALUE=19'b0000001_000000100010;
      15'b000_111110111110 : VALUE=19'b0000001_000000100001;
      15'b000_111110111111 : VALUE=19'b0000001_000000100001;
      15'b000_111111000000 : VALUE=19'b0000001_000000100000;
      15'b000_111111000001 : VALUE=19'b0000001_000000100000;
      15'b000_111111000010 : VALUE=19'b0000001_000000011111;
      15'b000_111111000011 : VALUE=19'b0000001_000000011111;
      15'b000_111111000100 : VALUE=19'b0000001_000000011110;
      15'b000_111111000101 : VALUE=19'b0000001_000000011110;
      15'b000_111111000110 : VALUE=19'b0000001_000000011101;
      15'b000_111111000111 : VALUE=19'b0000001_000000011101;
      15'b000_111111001000 : VALUE=19'b0000001_000000011100;
      15'b000_111111001001 : VALUE=19'b0000001_000000011100;
      15'b000_111111001010 : VALUE=19'b0000001_000000011011;
      15'b000_111111001011 : VALUE=19'b0000001_000000011011;
      15'b000_111111001100 : VALUE=19'b0000001_000000011010;
      15'b000_111111001101 : VALUE=19'b0000001_000000011010;
      15'b000_111111001110 : VALUE=19'b0000001_000000011001;
      15'b000_111111001111 : VALUE=19'b0000001_000000011001;
      15'b000_111111010000 : VALUE=19'b0000001_000000011000;
      15'b000_111111010001 : VALUE=19'b0000001_000000011000;
      15'b000_111111010010 : VALUE=19'b0000001_000000010111;
      15'b000_111111010011 : VALUE=19'b0000001_000000010111;
      15'b000_111111010100 : VALUE=19'b0000001_000000010110;
      15'b000_111111010101 : VALUE=19'b0000001_000000010110;
      15'b000_111111010110 : VALUE=19'b0000001_000000010101;
      15'b000_111111010111 : VALUE=19'b0000001_000000010101;
      15'b000_111111011000 : VALUE=19'b0000001_000000010100;
      15'b000_111111011001 : VALUE=19'b0000001_000000010100;
      15'b000_111111011010 : VALUE=19'b0000001_000000010011;
      15'b000_111111011011 : VALUE=19'b0000001_000000010011;
      15'b000_111111011100 : VALUE=19'b0000001_000000010010;
      15'b000_111111011101 : VALUE=19'b0000001_000000010010;
      15'b000_111111011110 : VALUE=19'b0000001_000000010001;
      15'b000_111111011111 : VALUE=19'b0000001_000000010001;
      15'b000_111111100000 : VALUE=19'b0000001_000000010000;
      15'b000_111111100001 : VALUE=19'b0000001_000000010000;
      15'b000_111111100010 : VALUE=19'b0000001_000000001111;
      15'b000_111111100011 : VALUE=19'b0000001_000000001111;
      15'b000_111111100100 : VALUE=19'b0000001_000000001110;
      15'b000_111111100101 : VALUE=19'b0000001_000000001110;
      15'b000_111111100110 : VALUE=19'b0000001_000000001101;
      15'b000_111111100111 : VALUE=19'b0000001_000000001101;
      15'b000_111111101000 : VALUE=19'b0000001_000000001100;
      15'b000_111111101001 : VALUE=19'b0000001_000000001100;
      15'b000_111111101010 : VALUE=19'b0000001_000000001011;
      15'b000_111111101011 : VALUE=19'b0000001_000000001011;
      15'b000_111111101100 : VALUE=19'b0000001_000000001010;
      15'b000_111111101101 : VALUE=19'b0000001_000000001010;
      15'b000_111111101110 : VALUE=19'b0000001_000000001001;
      15'b000_111111101111 : VALUE=19'b0000001_000000001001;
      15'b000_111111110000 : VALUE=19'b0000001_000000001000;
      15'b000_111111110001 : VALUE=19'b0000001_000000001000;
      15'b000_111111110010 : VALUE=19'b0000001_000000000111;
      15'b000_111111110011 : VALUE=19'b0000001_000000000111;
      15'b000_111111110100 : VALUE=19'b0000001_000000000110;
      15'b000_111111110101 : VALUE=19'b0000001_000000000110;
      15'b000_111111110110 : VALUE=19'b0000001_000000000101;
      15'b000_111111110111 : VALUE=19'b0000001_000000000101;
      15'b000_111111111000 : VALUE=19'b0000001_000000000100;
      15'b000_111111111001 : VALUE=19'b0000001_000000000100;
      15'b000_111111111010 : VALUE=19'b0000001_000000000011;
      15'b000_111111111011 : VALUE=19'b0000001_000000000011;
      15'b000_111111111100 : VALUE=19'b0000001_000000000010;
      15'b000_111111111101 : VALUE=19'b0000001_000000000010;
      15'b000_111111111110 : VALUE=19'b0000001_000000000001;
      15'b000_111111111111 : VALUE=19'b0000001_000000000001;
      15'b001_000000000000 : VALUE=19'b0000001_000000000000;
      15'b001_000000000001 : VALUE=19'b0000001_000000000000;
      15'b001_000000000010 : VALUE=19'b0000000_111111111111;
      15'b001_000000000011 : VALUE=19'b0000000_111111111111;
      15'b001_000000000100 : VALUE=19'b0000000_111111111110;
      15'b001_000000000101 : VALUE=19'b0000000_111111111110;
      15'b001_000000000110 : VALUE=19'b0000000_111111111101;
      15'b001_000000000111 : VALUE=19'b0000000_111111111101;
      15'b001_000000001000 : VALUE=19'b0000000_111111111100;
      15'b001_000000001001 : VALUE=19'b0000000_111111111100;
      15'b001_000000001010 : VALUE=19'b0000000_111111111011;
      15'b001_000000001011 : VALUE=19'b0000000_111111111011;
      15'b001_000000001100 : VALUE=19'b0000000_111111111010;
      15'b001_000000001101 : VALUE=19'b0000000_111111111010;
      15'b001_000000001110 : VALUE=19'b0000000_111111111001;
      15'b001_000000001111 : VALUE=19'b0000000_111111111001;
      15'b001_000000010000 : VALUE=19'b0000000_111111111000;
      15'b001_000000010001 : VALUE=19'b0000000_111111111000;
      15'b001_000000010010 : VALUE=19'b0000000_111111110111;
      15'b001_000000010011 : VALUE=19'b0000000_111111110111;
      15'b001_000000010100 : VALUE=19'b0000000_111111110110;
      15'b001_000000010101 : VALUE=19'b0000000_111111110110;
      15'b001_000000010110 : VALUE=19'b0000000_111111110101;
      15'b001_000000010111 : VALUE=19'b0000000_111111110101;
      15'b001_000000011000 : VALUE=19'b0000000_111111110100;
      15'b001_000000011001 : VALUE=19'b0000000_111111110100;
      15'b001_000000011010 : VALUE=19'b0000000_111111110011;
      15'b001_000000011011 : VALUE=19'b0000000_111111110011;
      15'b001_000000011100 : VALUE=19'b0000000_111111110010;
      15'b001_000000011101 : VALUE=19'b0000000_111111110010;
      15'b001_000000011110 : VALUE=19'b0000000_111111110001;
      15'b001_000000011111 : VALUE=19'b0000000_111111110001;
      15'b001_000000100000 : VALUE=19'b0000000_111111110000;
      15'b001_000000100001 : VALUE=19'b0000000_111111110000;
      15'b001_000000100010 : VALUE=19'b0000000_111111101111;
      15'b001_000000100011 : VALUE=19'b0000000_111111101111;
      15'b001_000000100100 : VALUE=19'b0000000_111111101110;
      15'b001_000000100101 : VALUE=19'b0000000_111111101110;
      15'b001_000000100110 : VALUE=19'b0000000_111111101101;
      15'b001_000000100111 : VALUE=19'b0000000_111111101101;
      15'b001_000000101000 : VALUE=19'b0000000_111111101100;
      15'b001_000000101001 : VALUE=19'b0000000_111111101100;
      15'b001_000000101010 : VALUE=19'b0000000_111111101011;
      15'b001_000000101011 : VALUE=19'b0000000_111111101011;
      15'b001_000000101100 : VALUE=19'b0000000_111111101010;
      15'b001_000000101101 : VALUE=19'b0000000_111111101010;
      15'b001_000000101110 : VALUE=19'b0000000_111111101001;
      15'b001_000000101111 : VALUE=19'b0000000_111111101001;
      15'b001_000000110000 : VALUE=19'b0000000_111111101000;
      15'b001_000000110001 : VALUE=19'b0000000_111111101000;
      15'b001_000000110010 : VALUE=19'b0000000_111111100111;
      15'b001_000000110011 : VALUE=19'b0000000_111111100111;
      15'b001_000000110100 : VALUE=19'b0000000_111111100110;
      15'b001_000000110101 : VALUE=19'b0000000_111111100110;
      15'b001_000000110110 : VALUE=19'b0000000_111111100101;
      15'b001_000000110111 : VALUE=19'b0000000_111111100101;
      15'b001_000000111000 : VALUE=19'b0000000_111111100100;
      15'b001_000000111001 : VALUE=19'b0000000_111111100100;
      15'b001_000000111010 : VALUE=19'b0000000_111111100011;
      15'b001_000000111011 : VALUE=19'b0000000_111111100011;
      15'b001_000000111100 : VALUE=19'b0000000_111111100010;
      15'b001_000000111101 : VALUE=19'b0000000_111111100010;
      15'b001_000000111110 : VALUE=19'b0000000_111111100001;
      15'b001_000000111111 : VALUE=19'b0000000_111111100001;
      15'b001_000001000000 : VALUE=19'b0000000_111111100000;
      15'b001_000001000001 : VALUE=19'b0000000_111111100000;
      15'b001_000001000010 : VALUE=19'b0000000_111111011111;
      15'b001_000001000011 : VALUE=19'b0000000_111111011111;
      15'b001_000001000100 : VALUE=19'b0000000_111111011110;
      15'b001_000001000101 : VALUE=19'b0000000_111111011110;
      15'b001_000001000110 : VALUE=19'b0000000_111111011101;
      15'b001_000001000111 : VALUE=19'b0000000_111111011101;
      15'b001_000001001000 : VALUE=19'b0000000_111111011100;
      15'b001_000001001001 : VALUE=19'b0000000_111111011100;
      15'b001_000001001010 : VALUE=19'b0000000_111111011011;
      15'b001_000001001011 : VALUE=19'b0000000_111111011011;
      15'b001_000001001100 : VALUE=19'b0000000_111111011011;
      15'b001_000001001101 : VALUE=19'b0000000_111111011010;
      15'b001_000001001110 : VALUE=19'b0000000_111111011010;
      15'b001_000001001111 : VALUE=19'b0000000_111111011001;
      15'b001_000001010000 : VALUE=19'b0000000_111111011001;
      15'b001_000001010001 : VALUE=19'b0000000_111111011000;
      15'b001_000001010010 : VALUE=19'b0000000_111111011000;
      15'b001_000001010011 : VALUE=19'b0000000_111111010111;
      15'b001_000001010100 : VALUE=19'b0000000_111111010111;
      15'b001_000001010101 : VALUE=19'b0000000_111111010110;
      15'b001_000001010110 : VALUE=19'b0000000_111111010110;
      15'b001_000001010111 : VALUE=19'b0000000_111111010101;
      15'b001_000001011000 : VALUE=19'b0000000_111111010101;
      15'b001_000001011001 : VALUE=19'b0000000_111111010100;
      15'b001_000001011010 : VALUE=19'b0000000_111111010100;
      15'b001_000001011011 : VALUE=19'b0000000_111111010011;
      15'b001_000001011100 : VALUE=19'b0000000_111111010011;
      15'b001_000001011101 : VALUE=19'b0000000_111111010010;
      15'b001_000001011110 : VALUE=19'b0000000_111111010010;
      15'b001_000001011111 : VALUE=19'b0000000_111111010001;
      15'b001_000001100000 : VALUE=19'b0000000_111111010001;
      15'b001_000001100001 : VALUE=19'b0000000_111111010000;
      15'b001_000001100010 : VALUE=19'b0000000_111111010000;
      15'b001_000001100011 : VALUE=19'b0000000_111111001111;
      15'b001_000001100100 : VALUE=19'b0000000_111111001111;
      15'b001_000001100101 : VALUE=19'b0000000_111111001110;
      15'b001_000001100110 : VALUE=19'b0000000_111111001110;
      15'b001_000001100111 : VALUE=19'b0000000_111111001101;
      15'b001_000001101000 : VALUE=19'b0000000_111111001101;
      15'b001_000001101001 : VALUE=19'b0000000_111111001100;
      15'b001_000001101010 : VALUE=19'b0000000_111111001100;
      15'b001_000001101011 : VALUE=19'b0000000_111111001100;
      15'b001_000001101100 : VALUE=19'b0000000_111111001011;
      15'b001_000001101101 : VALUE=19'b0000000_111111001011;
      15'b001_000001101110 : VALUE=19'b0000000_111111001010;
      15'b001_000001101111 : VALUE=19'b0000000_111111001010;
      15'b001_000001110000 : VALUE=19'b0000000_111111001001;
      15'b001_000001110001 : VALUE=19'b0000000_111111001001;
      15'b001_000001110010 : VALUE=19'b0000000_111111001000;
      15'b001_000001110011 : VALUE=19'b0000000_111111001000;
      15'b001_000001110100 : VALUE=19'b0000000_111111000111;
      15'b001_000001110101 : VALUE=19'b0000000_111111000111;
      15'b001_000001110110 : VALUE=19'b0000000_111111000110;
      15'b001_000001110111 : VALUE=19'b0000000_111111000110;
      15'b001_000001111000 : VALUE=19'b0000000_111111000101;
      15'b001_000001111001 : VALUE=19'b0000000_111111000101;
      15'b001_000001111010 : VALUE=19'b0000000_111111000100;
      15'b001_000001111011 : VALUE=19'b0000000_111111000100;
      15'b001_000001111100 : VALUE=19'b0000000_111111000011;
      15'b001_000001111101 : VALUE=19'b0000000_111111000011;
      15'b001_000001111110 : VALUE=19'b0000000_111111000010;
      15'b001_000001111111 : VALUE=19'b0000000_111111000010;
      15'b001_000010000000 : VALUE=19'b0000000_111111000001;
      15'b001_000010000001 : VALUE=19'b0000000_111111000001;
      15'b001_000010000010 : VALUE=19'b0000000_111111000001;
      15'b001_000010000011 : VALUE=19'b0000000_111111000000;
      15'b001_000010000100 : VALUE=19'b0000000_111111000000;
      15'b001_000010000101 : VALUE=19'b0000000_111110111111;
      15'b001_000010000110 : VALUE=19'b0000000_111110111111;
      15'b001_000010000111 : VALUE=19'b0000000_111110111110;
      15'b001_000010001000 : VALUE=19'b0000000_111110111110;
      15'b001_000010001001 : VALUE=19'b0000000_111110111101;
      15'b001_000010001010 : VALUE=19'b0000000_111110111101;
      15'b001_000010001011 : VALUE=19'b0000000_111110111100;
      15'b001_000010001100 : VALUE=19'b0000000_111110111100;
      15'b001_000010001101 : VALUE=19'b0000000_111110111011;
      15'b001_000010001110 : VALUE=19'b0000000_111110111011;
      15'b001_000010001111 : VALUE=19'b0000000_111110111010;
      15'b001_000010010000 : VALUE=19'b0000000_111110111010;
      15'b001_000010010001 : VALUE=19'b0000000_111110111001;
      15'b001_000010010010 : VALUE=19'b0000000_111110111001;
      15'b001_000010010011 : VALUE=19'b0000000_111110111000;
      15'b001_000010010100 : VALUE=19'b0000000_111110111000;
      15'b001_000010010101 : VALUE=19'b0000000_111110110111;
      15'b001_000010010110 : VALUE=19'b0000000_111110110111;
      15'b001_000010010111 : VALUE=19'b0000000_111110110111;
      15'b001_000010011000 : VALUE=19'b0000000_111110110110;
      15'b001_000010011001 : VALUE=19'b0000000_111110110110;
      15'b001_000010011010 : VALUE=19'b0000000_111110110101;
      15'b001_000010011011 : VALUE=19'b0000000_111110110101;
      15'b001_000010011100 : VALUE=19'b0000000_111110110100;
      15'b001_000010011101 : VALUE=19'b0000000_111110110100;
      15'b001_000010011110 : VALUE=19'b0000000_111110110011;
      15'b001_000010011111 : VALUE=19'b0000000_111110110011;
      15'b001_000010100000 : VALUE=19'b0000000_111110110010;
      15'b001_000010100001 : VALUE=19'b0000000_111110110010;
      15'b001_000010100010 : VALUE=19'b0000000_111110110001;
      15'b001_000010100011 : VALUE=19'b0000000_111110110001;
      15'b001_000010100100 : VALUE=19'b0000000_111110110000;
      15'b001_000010100101 : VALUE=19'b0000000_111110110000;
      15'b001_000010100110 : VALUE=19'b0000000_111110101111;
      15'b001_000010100111 : VALUE=19'b0000000_111110101111;
      15'b001_000010101000 : VALUE=19'b0000000_111110101110;
      15'b001_000010101001 : VALUE=19'b0000000_111110101110;
      15'b001_000010101010 : VALUE=19'b0000000_111110101110;
      15'b001_000010101011 : VALUE=19'b0000000_111110101101;
      15'b001_000010101100 : VALUE=19'b0000000_111110101101;
      15'b001_000010101101 : VALUE=19'b0000000_111110101100;
      15'b001_000010101110 : VALUE=19'b0000000_111110101100;
      15'b001_000010101111 : VALUE=19'b0000000_111110101011;
      15'b001_000010110000 : VALUE=19'b0000000_111110101011;
      15'b001_000010110001 : VALUE=19'b0000000_111110101010;
      15'b001_000010110010 : VALUE=19'b0000000_111110101010;
      15'b001_000010110011 : VALUE=19'b0000000_111110101001;
      15'b001_000010110100 : VALUE=19'b0000000_111110101001;
      15'b001_000010110101 : VALUE=19'b0000000_111110101000;
      15'b001_000010110110 : VALUE=19'b0000000_111110101000;
      15'b001_000010110111 : VALUE=19'b0000000_111110100111;
      15'b001_000010111000 : VALUE=19'b0000000_111110100111;
      15'b001_000010111001 : VALUE=19'b0000000_111110100111;
      15'b001_000010111010 : VALUE=19'b0000000_111110100110;
      15'b001_000010111011 : VALUE=19'b0000000_111110100110;
      15'b001_000010111100 : VALUE=19'b0000000_111110100101;
      15'b001_000010111101 : VALUE=19'b0000000_111110100101;
      15'b001_000010111110 : VALUE=19'b0000000_111110100100;
      15'b001_000010111111 : VALUE=19'b0000000_111110100100;
      15'b001_000011000000 : VALUE=19'b0000000_111110100011;
      15'b001_000011000001 : VALUE=19'b0000000_111110100011;
      15'b001_000011000010 : VALUE=19'b0000000_111110100010;
      15'b001_000011000011 : VALUE=19'b0000000_111110100010;
      15'b001_000011000100 : VALUE=19'b0000000_111110100001;
      15'b001_000011000101 : VALUE=19'b0000000_111110100001;
      15'b001_000011000110 : VALUE=19'b0000000_111110100000;
      15'b001_000011000111 : VALUE=19'b0000000_111110100000;
      15'b001_000011001000 : VALUE=19'b0000000_111110100000;
      15'b001_000011001001 : VALUE=19'b0000000_111110011111;
      15'b001_000011001010 : VALUE=19'b0000000_111110011111;
      15'b001_000011001011 : VALUE=19'b0000000_111110011110;
      15'b001_000011001100 : VALUE=19'b0000000_111110011110;
      15'b001_000011001101 : VALUE=19'b0000000_111110011101;
      15'b001_000011001110 : VALUE=19'b0000000_111110011101;
      15'b001_000011001111 : VALUE=19'b0000000_111110011100;
      15'b001_000011010000 : VALUE=19'b0000000_111110011100;
      15'b001_000011010001 : VALUE=19'b0000000_111110011011;
      15'b001_000011010010 : VALUE=19'b0000000_111110011011;
      15'b001_000011010011 : VALUE=19'b0000000_111110011010;
      15'b001_000011010100 : VALUE=19'b0000000_111110011010;
      15'b001_000011010101 : VALUE=19'b0000000_111110011001;
      15'b001_000011010110 : VALUE=19'b0000000_111110011001;
      15'b001_000011010111 : VALUE=19'b0000000_111110011001;
      15'b001_000011011000 : VALUE=19'b0000000_111110011000;
      15'b001_000011011001 : VALUE=19'b0000000_111110011000;
      15'b001_000011011010 : VALUE=19'b0000000_111110010111;
      15'b001_000011011011 : VALUE=19'b0000000_111110010111;
      15'b001_000011011100 : VALUE=19'b0000000_111110010110;
      15'b001_000011011101 : VALUE=19'b0000000_111110010110;
      15'b001_000011011110 : VALUE=19'b0000000_111110010101;
      15'b001_000011011111 : VALUE=19'b0000000_111110010101;
      15'b001_000011100000 : VALUE=19'b0000000_111110010100;
      15'b001_000011100001 : VALUE=19'b0000000_111110010100;
      15'b001_000011100010 : VALUE=19'b0000000_111110010011;
      15'b001_000011100011 : VALUE=19'b0000000_111110010011;
      15'b001_000011100100 : VALUE=19'b0000000_111110010011;
      15'b001_000011100101 : VALUE=19'b0000000_111110010010;
      15'b001_000011100110 : VALUE=19'b0000000_111110010010;
      15'b001_000011100111 : VALUE=19'b0000000_111110010001;
      15'b001_000011101000 : VALUE=19'b0000000_111110010001;
      15'b001_000011101001 : VALUE=19'b0000000_111110010000;
      15'b001_000011101010 : VALUE=19'b0000000_111110010000;
      15'b001_000011101011 : VALUE=19'b0000000_111110001111;
      15'b001_000011101100 : VALUE=19'b0000000_111110001111;
      15'b001_000011101101 : VALUE=19'b0000000_111110001110;
      15'b001_000011101110 : VALUE=19'b0000000_111110001110;
      15'b001_000011101111 : VALUE=19'b0000000_111110001101;
      15'b001_000011110000 : VALUE=19'b0000000_111110001101;
      15'b001_000011110001 : VALUE=19'b0000000_111110001101;
      15'b001_000011110010 : VALUE=19'b0000000_111110001100;
      15'b001_000011110011 : VALUE=19'b0000000_111110001100;
      15'b001_000011110100 : VALUE=19'b0000000_111110001011;
      15'b001_000011110101 : VALUE=19'b0000000_111110001011;
      15'b001_000011110110 : VALUE=19'b0000000_111110001010;
      15'b001_000011110111 : VALUE=19'b0000000_111110001010;
      15'b001_000011111000 : VALUE=19'b0000000_111110001001;
      15'b001_000011111001 : VALUE=19'b0000000_111110001001;
      15'b001_000011111010 : VALUE=19'b0000000_111110001000;
      15'b001_000011111011 : VALUE=19'b0000000_111110001000;
      15'b001_000011111100 : VALUE=19'b0000000_111110001000;
      15'b001_000011111101 : VALUE=19'b0000000_111110000111;
      15'b001_000011111110 : VALUE=19'b0000000_111110000111;
      15'b001_000011111111 : VALUE=19'b0000000_111110000110;
      15'b001_000100000000 : VALUE=19'b0000000_111110000110;
      15'b001_000100000001 : VALUE=19'b0000000_111110000101;
      15'b001_000100000010 : VALUE=19'b0000000_111110000101;
      15'b001_000100000011 : VALUE=19'b0000000_111110000100;
      15'b001_000100000100 : VALUE=19'b0000000_111110000100;
      15'b001_000100000101 : VALUE=19'b0000000_111110000011;
      15'b001_000100000110 : VALUE=19'b0000000_111110000011;
      15'b001_000100000111 : VALUE=19'b0000000_111110000011;
      15'b001_000100001000 : VALUE=19'b0000000_111110000010;
      15'b001_000100001001 : VALUE=19'b0000000_111110000010;
      15'b001_000100001010 : VALUE=19'b0000000_111110000001;
      15'b001_000100001011 : VALUE=19'b0000000_111110000001;
      15'b001_000100001100 : VALUE=19'b0000000_111110000000;
      15'b001_000100001101 : VALUE=19'b0000000_111110000000;
      15'b001_000100001110 : VALUE=19'b0000000_111101111111;
      15'b001_000100001111 : VALUE=19'b0000000_111101111111;
      15'b001_000100010000 : VALUE=19'b0000000_111101111110;
      15'b001_000100010001 : VALUE=19'b0000000_111101111110;
      15'b001_000100010010 : VALUE=19'b0000000_111101111110;
      15'b001_000100010011 : VALUE=19'b0000000_111101111101;
      15'b001_000100010100 : VALUE=19'b0000000_111101111101;
      15'b001_000100010101 : VALUE=19'b0000000_111101111100;
      15'b001_000100010110 : VALUE=19'b0000000_111101111100;
      15'b001_000100010111 : VALUE=19'b0000000_111101111011;
      15'b001_000100011000 : VALUE=19'b0000000_111101111011;
      15'b001_000100011001 : VALUE=19'b0000000_111101111010;
      15'b001_000100011010 : VALUE=19'b0000000_111101111010;
      15'b001_000100011011 : VALUE=19'b0000000_111101111001;
      15'b001_000100011100 : VALUE=19'b0000000_111101111001;
      15'b001_000100011101 : VALUE=19'b0000000_111101111001;
      15'b001_000100011110 : VALUE=19'b0000000_111101111000;
      15'b001_000100011111 : VALUE=19'b0000000_111101111000;
      15'b001_000100100000 : VALUE=19'b0000000_111101110111;
      15'b001_000100100001 : VALUE=19'b0000000_111101110111;
      15'b001_000100100010 : VALUE=19'b0000000_111101110110;
      15'b001_000100100011 : VALUE=19'b0000000_111101110110;
      15'b001_000100100100 : VALUE=19'b0000000_111101110101;
      15'b001_000100100101 : VALUE=19'b0000000_111101110101;
      15'b001_000100100110 : VALUE=19'b0000000_111101110100;
      15'b001_000100100111 : VALUE=19'b0000000_111101110100;
      15'b001_000100101000 : VALUE=19'b0000000_111101110100;
      15'b001_000100101001 : VALUE=19'b0000000_111101110011;
      15'b001_000100101010 : VALUE=19'b0000000_111101110011;
      15'b001_000100101011 : VALUE=19'b0000000_111101110010;
      15'b001_000100101100 : VALUE=19'b0000000_111101110010;
      15'b001_000100101101 : VALUE=19'b0000000_111101110001;
      15'b001_000100101110 : VALUE=19'b0000000_111101110001;
      15'b001_000100101111 : VALUE=19'b0000000_111101110000;
      15'b001_000100110000 : VALUE=19'b0000000_111101110000;
      15'b001_000100110001 : VALUE=19'b0000000_111101110000;
      15'b001_000100110010 : VALUE=19'b0000000_111101101111;
      15'b001_000100110011 : VALUE=19'b0000000_111101101111;
      15'b001_000100110100 : VALUE=19'b0000000_111101101110;
      15'b001_000100110101 : VALUE=19'b0000000_111101101110;
      15'b001_000100110110 : VALUE=19'b0000000_111101101101;
      15'b001_000100110111 : VALUE=19'b0000000_111101101101;
      15'b001_000100111000 : VALUE=19'b0000000_111101101100;
      15'b001_000100111001 : VALUE=19'b0000000_111101101100;
      15'b001_000100111010 : VALUE=19'b0000000_111101101011;
      15'b001_000100111011 : VALUE=19'b0000000_111101101011;
      15'b001_000100111100 : VALUE=19'b0000000_111101101011;
      15'b001_000100111101 : VALUE=19'b0000000_111101101010;
      15'b001_000100111110 : VALUE=19'b0000000_111101101010;
      15'b001_000100111111 : VALUE=19'b0000000_111101101001;
      15'b001_000101000000 : VALUE=19'b0000000_111101101001;
      15'b001_000101000001 : VALUE=19'b0000000_111101101000;
      15'b001_000101000010 : VALUE=19'b0000000_111101101000;
      15'b001_000101000011 : VALUE=19'b0000000_111101100111;
      15'b001_000101000100 : VALUE=19'b0000000_111101100111;
      15'b001_000101000101 : VALUE=19'b0000000_111101100111;
      15'b001_000101000110 : VALUE=19'b0000000_111101100110;
      15'b001_000101000111 : VALUE=19'b0000000_111101100110;
      15'b001_000101001000 : VALUE=19'b0000000_111101100101;
      15'b001_000101001001 : VALUE=19'b0000000_111101100101;
      15'b001_000101001010 : VALUE=19'b0000000_111101100100;
      15'b001_000101001011 : VALUE=19'b0000000_111101100100;
      15'b001_000101001100 : VALUE=19'b0000000_111101100011;
      15'b001_000101001101 : VALUE=19'b0000000_111101100011;
      15'b001_000101001110 : VALUE=19'b0000000_111101100011;
      15'b001_000101001111 : VALUE=19'b0000000_111101100010;
      15'b001_000101010000 : VALUE=19'b0000000_111101100010;
      15'b001_000101010001 : VALUE=19'b0000000_111101100001;
      15'b001_000101010010 : VALUE=19'b0000000_111101100001;
      15'b001_000101010011 : VALUE=19'b0000000_111101100000;
      15'b001_000101010100 : VALUE=19'b0000000_111101100000;
      15'b001_000101010101 : VALUE=19'b0000000_111101011111;
      15'b001_000101010110 : VALUE=19'b0000000_111101011111;
      15'b001_000101010111 : VALUE=19'b0000000_111101011111;
      15'b001_000101011000 : VALUE=19'b0000000_111101011110;
      15'b001_000101011001 : VALUE=19'b0000000_111101011110;
      15'b001_000101011010 : VALUE=19'b0000000_111101011101;
      15'b001_000101011011 : VALUE=19'b0000000_111101011101;
      15'b001_000101011100 : VALUE=19'b0000000_111101011100;
      15'b001_000101011101 : VALUE=19'b0000000_111101011100;
      15'b001_000101011110 : VALUE=19'b0000000_111101011011;
      15'b001_000101011111 : VALUE=19'b0000000_111101011011;
      15'b001_000101100000 : VALUE=19'b0000000_111101011011;
      15'b001_000101100001 : VALUE=19'b0000000_111101011010;
      15'b001_000101100010 : VALUE=19'b0000000_111101011010;
      15'b001_000101100011 : VALUE=19'b0000000_111101011001;
      15'b001_000101100100 : VALUE=19'b0000000_111101011001;
      15'b001_000101100101 : VALUE=19'b0000000_111101011000;
      15'b001_000101100110 : VALUE=19'b0000000_111101011000;
      15'b001_000101100111 : VALUE=19'b0000000_111101010111;
      15'b001_000101101000 : VALUE=19'b0000000_111101010111;
      15'b001_000101101001 : VALUE=19'b0000000_111101010111;
      15'b001_000101101010 : VALUE=19'b0000000_111101010110;
      15'b001_000101101011 : VALUE=19'b0000000_111101010110;
      15'b001_000101101100 : VALUE=19'b0000000_111101010101;
      15'b001_000101101101 : VALUE=19'b0000000_111101010101;
      15'b001_000101101110 : VALUE=19'b0000000_111101010100;
      15'b001_000101101111 : VALUE=19'b0000000_111101010100;
      15'b001_000101110000 : VALUE=19'b0000000_111101010100;
      15'b001_000101110001 : VALUE=19'b0000000_111101010011;
      15'b001_000101110010 : VALUE=19'b0000000_111101010011;
      15'b001_000101110011 : VALUE=19'b0000000_111101010010;
      15'b001_000101110100 : VALUE=19'b0000000_111101010010;
      15'b001_000101110101 : VALUE=19'b0000000_111101010001;
      15'b001_000101110110 : VALUE=19'b0000000_111101010001;
      15'b001_000101110111 : VALUE=19'b0000000_111101010000;
      15'b001_000101111000 : VALUE=19'b0000000_111101010000;
      15'b001_000101111001 : VALUE=19'b0000000_111101010000;
      15'b001_000101111010 : VALUE=19'b0000000_111101001111;
      15'b001_000101111011 : VALUE=19'b0000000_111101001111;
      15'b001_000101111100 : VALUE=19'b0000000_111101001110;
      15'b001_000101111101 : VALUE=19'b0000000_111101001110;
      15'b001_000101111110 : VALUE=19'b0000000_111101001101;
      15'b001_000101111111 : VALUE=19'b0000000_111101001101;
      15'b001_000110000000 : VALUE=19'b0000000_111101001101;
      15'b001_000110000001 : VALUE=19'b0000000_111101001100;
      15'b001_000110000010 : VALUE=19'b0000000_111101001100;
      15'b001_000110000011 : VALUE=19'b0000000_111101001011;
      15'b001_000110000100 : VALUE=19'b0000000_111101001011;
      15'b001_000110000101 : VALUE=19'b0000000_111101001010;
      15'b001_000110000110 : VALUE=19'b0000000_111101001010;
      15'b001_000110000111 : VALUE=19'b0000000_111101001001;
      15'b001_000110001000 : VALUE=19'b0000000_111101001001;
      15'b001_000110001001 : VALUE=19'b0000000_111101001001;
      15'b001_000110001010 : VALUE=19'b0000000_111101001000;
      15'b001_000110001011 : VALUE=19'b0000000_111101001000;
      15'b001_000110001100 : VALUE=19'b0000000_111101000111;
      15'b001_000110001101 : VALUE=19'b0000000_111101000111;
      15'b001_000110001110 : VALUE=19'b0000000_111101000110;
      15'b001_000110001111 : VALUE=19'b0000000_111101000110;
      15'b001_000110010000 : VALUE=19'b0000000_111101000110;
      15'b001_000110010001 : VALUE=19'b0000000_111101000101;
      15'b001_000110010010 : VALUE=19'b0000000_111101000101;
      15'b001_000110010011 : VALUE=19'b0000000_111101000100;
      15'b001_000110010100 : VALUE=19'b0000000_111101000100;
      15'b001_000110010101 : VALUE=19'b0000000_111101000011;
      15'b001_000110010110 : VALUE=19'b0000000_111101000011;
      15'b001_000110010111 : VALUE=19'b0000000_111101000011;
      15'b001_000110011000 : VALUE=19'b0000000_111101000010;
      15'b001_000110011001 : VALUE=19'b0000000_111101000010;
      15'b001_000110011010 : VALUE=19'b0000000_111101000001;
      15'b001_000110011011 : VALUE=19'b0000000_111101000001;
      15'b001_000110011100 : VALUE=19'b0000000_111101000000;
      15'b001_000110011101 : VALUE=19'b0000000_111101000000;
      15'b001_000110011110 : VALUE=19'b0000000_111100111111;
      15'b001_000110011111 : VALUE=19'b0000000_111100111111;
      15'b001_000110100000 : VALUE=19'b0000000_111100111111;
      15'b001_000110100001 : VALUE=19'b0000000_111100111110;
      15'b001_000110100010 : VALUE=19'b0000000_111100111110;
      15'b001_000110100011 : VALUE=19'b0000000_111100111101;
      15'b001_000110100100 : VALUE=19'b0000000_111100111101;
      15'b001_000110100101 : VALUE=19'b0000000_111100111100;
      15'b001_000110100110 : VALUE=19'b0000000_111100111100;
      15'b001_000110100111 : VALUE=19'b0000000_111100111100;
      15'b001_000110101000 : VALUE=19'b0000000_111100111011;
      15'b001_000110101001 : VALUE=19'b0000000_111100111011;
      15'b001_000110101010 : VALUE=19'b0000000_111100111010;
      15'b001_000110101011 : VALUE=19'b0000000_111100111010;
      15'b001_000110101100 : VALUE=19'b0000000_111100111001;
      15'b001_000110101101 : VALUE=19'b0000000_111100111001;
      15'b001_000110101110 : VALUE=19'b0000000_111100111001;
      15'b001_000110101111 : VALUE=19'b0000000_111100111000;
      15'b001_000110110000 : VALUE=19'b0000000_111100111000;
      15'b001_000110110001 : VALUE=19'b0000000_111100110111;
      15'b001_000110110010 : VALUE=19'b0000000_111100110111;
      15'b001_000110110011 : VALUE=19'b0000000_111100110110;
      15'b001_000110110100 : VALUE=19'b0000000_111100110110;
      15'b001_000110110101 : VALUE=19'b0000000_111100110110;
      15'b001_000110110110 : VALUE=19'b0000000_111100110101;
      15'b001_000110110111 : VALUE=19'b0000000_111100110101;
      15'b001_000110111000 : VALUE=19'b0000000_111100110100;
      15'b001_000110111001 : VALUE=19'b0000000_111100110100;
      15'b001_000110111010 : VALUE=19'b0000000_111100110011;
      15'b001_000110111011 : VALUE=19'b0000000_111100110011;
      15'b001_000110111100 : VALUE=19'b0000000_111100110011;
      15'b001_000110111101 : VALUE=19'b0000000_111100110010;
      15'b001_000110111110 : VALUE=19'b0000000_111100110010;
      15'b001_000110111111 : VALUE=19'b0000000_111100110001;
      15'b001_000111000000 : VALUE=19'b0000000_111100110001;
      15'b001_000111000001 : VALUE=19'b0000000_111100110000;
      15'b001_000111000010 : VALUE=19'b0000000_111100110000;
      15'b001_000111000011 : VALUE=19'b0000000_111100110000;
      15'b001_000111000100 : VALUE=19'b0000000_111100101111;
      15'b001_000111000101 : VALUE=19'b0000000_111100101111;
      15'b001_000111000110 : VALUE=19'b0000000_111100101110;
      15'b001_000111000111 : VALUE=19'b0000000_111100101110;
      15'b001_000111001000 : VALUE=19'b0000000_111100101101;
      15'b001_000111001001 : VALUE=19'b0000000_111100101101;
      15'b001_000111001010 : VALUE=19'b0000000_111100101101;
      15'b001_000111001011 : VALUE=19'b0000000_111100101100;
      15'b001_000111001100 : VALUE=19'b0000000_111100101100;
      15'b001_000111001101 : VALUE=19'b0000000_111100101011;
      15'b001_000111001110 : VALUE=19'b0000000_111100101011;
      15'b001_000111001111 : VALUE=19'b0000000_111100101010;
      15'b001_000111010000 : VALUE=19'b0000000_111100101010;
      15'b001_000111010001 : VALUE=19'b0000000_111100101010;
      15'b001_000111010010 : VALUE=19'b0000000_111100101001;
      15'b001_000111010011 : VALUE=19'b0000000_111100101001;
      15'b001_000111010100 : VALUE=19'b0000000_111100101000;
      15'b001_000111010101 : VALUE=19'b0000000_111100101000;
      15'b001_000111010110 : VALUE=19'b0000000_111100100111;
      15'b001_000111010111 : VALUE=19'b0000000_111100100111;
      15'b001_000111011000 : VALUE=19'b0000000_111100100111;
      15'b001_000111011001 : VALUE=19'b0000000_111100100110;
      15'b001_000111011010 : VALUE=19'b0000000_111100100110;
      15'b001_000111011011 : VALUE=19'b0000000_111100100101;
      15'b001_000111011100 : VALUE=19'b0000000_111100100101;
      15'b001_000111011101 : VALUE=19'b0000000_111100100100;
      15'b001_000111011110 : VALUE=19'b0000000_111100100100;
      15'b001_000111011111 : VALUE=19'b0000000_111100100100;
      15'b001_000111100000 : VALUE=19'b0000000_111100100011;
      15'b001_000111100001 : VALUE=19'b0000000_111100100011;
      15'b001_000111100010 : VALUE=19'b0000000_111100100010;
      15'b001_000111100011 : VALUE=19'b0000000_111100100010;
      15'b001_000111100100 : VALUE=19'b0000000_111100100010;
      15'b001_000111100101 : VALUE=19'b0000000_111100100001;
      15'b001_000111100110 : VALUE=19'b0000000_111100100001;
      15'b001_000111100111 : VALUE=19'b0000000_111100100000;
      15'b001_000111101000 : VALUE=19'b0000000_111100100000;
      15'b001_000111101001 : VALUE=19'b0000000_111100011111;
      15'b001_000111101010 : VALUE=19'b0000000_111100011111;
      15'b001_000111101011 : VALUE=19'b0000000_111100011111;
      15'b001_000111101100 : VALUE=19'b0000000_111100011110;
      15'b001_000111101101 : VALUE=19'b0000000_111100011110;
      15'b001_000111101110 : VALUE=19'b0000000_111100011101;
      15'b001_000111101111 : VALUE=19'b0000000_111100011101;
      15'b001_000111110000 : VALUE=19'b0000000_111100011100;
      15'b001_000111110001 : VALUE=19'b0000000_111100011100;
      15'b001_000111110010 : VALUE=19'b0000000_111100011100;
      15'b001_000111110011 : VALUE=19'b0000000_111100011011;
      15'b001_000111110100 : VALUE=19'b0000000_111100011011;
      15'b001_000111110101 : VALUE=19'b0000000_111100011010;
      15'b001_000111110110 : VALUE=19'b0000000_111100011010;
      15'b001_000111110111 : VALUE=19'b0000000_111100011010;
      15'b001_000111111000 : VALUE=19'b0000000_111100011001;
      15'b001_000111111001 : VALUE=19'b0000000_111100011001;
      15'b001_000111111010 : VALUE=19'b0000000_111100011000;
      15'b001_000111111011 : VALUE=19'b0000000_111100011000;
      15'b001_000111111100 : VALUE=19'b0000000_111100010111;
      15'b001_000111111101 : VALUE=19'b0000000_111100010111;
      15'b001_000111111110 : VALUE=19'b0000000_111100010111;
      15'b001_000111111111 : VALUE=19'b0000000_111100010110;
      15'b001_001000000000 : VALUE=19'b0000000_111100010110;
      15'b001_001000000001 : VALUE=19'b0000000_111100010101;
      15'b001_001000000010 : VALUE=19'b0000000_111100010101;
      15'b001_001000000011 : VALUE=19'b0000000_111100010100;
      15'b001_001000000100 : VALUE=19'b0000000_111100010100;
      15'b001_001000000101 : VALUE=19'b0000000_111100010100;
      15'b001_001000000110 : VALUE=19'b0000000_111100010011;
      15'b001_001000000111 : VALUE=19'b0000000_111100010011;
      15'b001_001000001000 : VALUE=19'b0000000_111100010010;
      15'b001_001000001001 : VALUE=19'b0000000_111100010010;
      15'b001_001000001010 : VALUE=19'b0000000_111100010010;
      15'b001_001000001011 : VALUE=19'b0000000_111100010001;
      15'b001_001000001100 : VALUE=19'b0000000_111100010001;
      15'b001_001000001101 : VALUE=19'b0000000_111100010000;
      15'b001_001000001110 : VALUE=19'b0000000_111100010000;
      15'b001_001000001111 : VALUE=19'b0000000_111100001111;
      15'b001_001000010000 : VALUE=19'b0000000_111100001111;
      15'b001_001000010001 : VALUE=19'b0000000_111100001111;
      15'b001_001000010010 : VALUE=19'b0000000_111100001110;
      15'b001_001000010011 : VALUE=19'b0000000_111100001110;
      15'b001_001000010100 : VALUE=19'b0000000_111100001101;
      15'b001_001000010101 : VALUE=19'b0000000_111100001101;
      15'b001_001000010110 : VALUE=19'b0000000_111100001101;
      15'b001_001000010111 : VALUE=19'b0000000_111100001100;
      15'b001_001000011000 : VALUE=19'b0000000_111100001100;
      15'b001_001000011001 : VALUE=19'b0000000_111100001011;
      15'b001_001000011010 : VALUE=19'b0000000_111100001011;
      15'b001_001000011011 : VALUE=19'b0000000_111100001010;
      15'b001_001000011100 : VALUE=19'b0000000_111100001010;
      15'b001_001000011101 : VALUE=19'b0000000_111100001010;
      15'b001_001000011110 : VALUE=19'b0000000_111100001001;
      15'b001_001000011111 : VALUE=19'b0000000_111100001001;
      15'b001_001000100000 : VALUE=19'b0000000_111100001000;
      15'b001_001000100001 : VALUE=19'b0000000_111100001000;
      15'b001_001000100010 : VALUE=19'b0000000_111100001000;
      15'b001_001000100011 : VALUE=19'b0000000_111100000111;
      15'b001_001000100100 : VALUE=19'b0000000_111100000111;
      15'b001_001000100101 : VALUE=19'b0000000_111100000110;
      15'b001_001000100110 : VALUE=19'b0000000_111100000110;
      15'b001_001000100111 : VALUE=19'b0000000_111100000110;
      15'b001_001000101000 : VALUE=19'b0000000_111100000101;
      15'b001_001000101001 : VALUE=19'b0000000_111100000101;
      15'b001_001000101010 : VALUE=19'b0000000_111100000100;
      15'b001_001000101011 : VALUE=19'b0000000_111100000100;
      15'b001_001000101100 : VALUE=19'b0000000_111100000011;
      15'b001_001000101101 : VALUE=19'b0000000_111100000011;
      15'b001_001000101110 : VALUE=19'b0000000_111100000011;
      15'b001_001000101111 : VALUE=19'b0000000_111100000010;
      15'b001_001000110000 : VALUE=19'b0000000_111100000010;
      15'b001_001000110001 : VALUE=19'b0000000_111100000001;
      15'b001_001000110010 : VALUE=19'b0000000_111100000001;
      15'b001_001000110011 : VALUE=19'b0000000_111100000001;
      15'b001_001000110100 : VALUE=19'b0000000_111100000000;
      15'b001_001000110101 : VALUE=19'b0000000_111100000000;
      15'b001_001000110110 : VALUE=19'b0000000_111011111111;
      15'b001_001000110111 : VALUE=19'b0000000_111011111111;
      15'b001_001000111000 : VALUE=19'b0000000_111011111110;
      15'b001_001000111001 : VALUE=19'b0000000_111011111110;
      15'b001_001000111010 : VALUE=19'b0000000_111011111110;
      15'b001_001000111011 : VALUE=19'b0000000_111011111101;
      15'b001_001000111100 : VALUE=19'b0000000_111011111101;
      15'b001_001000111101 : VALUE=19'b0000000_111011111100;
      15'b001_001000111110 : VALUE=19'b0000000_111011111100;
      15'b001_001000111111 : VALUE=19'b0000000_111011111100;
      15'b001_001001000000 : VALUE=19'b0000000_111011111011;
      15'b001_001001000001 : VALUE=19'b0000000_111011111011;
      15'b001_001001000010 : VALUE=19'b0000000_111011111010;
      15'b001_001001000011 : VALUE=19'b0000000_111011111010;
      15'b001_001001000100 : VALUE=19'b0000000_111011111010;
      15'b001_001001000101 : VALUE=19'b0000000_111011111001;
      15'b001_001001000110 : VALUE=19'b0000000_111011111001;
      15'b001_001001000111 : VALUE=19'b0000000_111011111000;
      15'b001_001001001000 : VALUE=19'b0000000_111011111000;
      15'b001_001001001001 : VALUE=19'b0000000_111011111000;
      15'b001_001001001010 : VALUE=19'b0000000_111011110111;
      15'b001_001001001011 : VALUE=19'b0000000_111011110111;
      15'b001_001001001100 : VALUE=19'b0000000_111011110110;
      15'b001_001001001101 : VALUE=19'b0000000_111011110110;
      15'b001_001001001110 : VALUE=19'b0000000_111011110101;
      15'b001_001001001111 : VALUE=19'b0000000_111011110101;
      15'b001_001001010000 : VALUE=19'b0000000_111011110101;
      15'b001_001001010001 : VALUE=19'b0000000_111011110100;
      15'b001_001001010010 : VALUE=19'b0000000_111011110100;
      15'b001_001001010011 : VALUE=19'b0000000_111011110011;
      15'b001_001001010100 : VALUE=19'b0000000_111011110011;
      15'b001_001001010101 : VALUE=19'b0000000_111011110011;
      15'b001_001001010110 : VALUE=19'b0000000_111011110010;
      15'b001_001001010111 : VALUE=19'b0000000_111011110010;
      15'b001_001001011000 : VALUE=19'b0000000_111011110001;
      15'b001_001001011001 : VALUE=19'b0000000_111011110001;
      15'b001_001001011010 : VALUE=19'b0000000_111011110001;
      15'b001_001001011011 : VALUE=19'b0000000_111011110000;
      15'b001_001001011100 : VALUE=19'b0000000_111011110000;
      15'b001_001001011101 : VALUE=19'b0000000_111011101111;
      15'b001_001001011110 : VALUE=19'b0000000_111011101111;
      15'b001_001001011111 : VALUE=19'b0000000_111011101111;
      15'b001_001001100000 : VALUE=19'b0000000_111011101110;
      15'b001_001001100001 : VALUE=19'b0000000_111011101110;
      15'b001_001001100010 : VALUE=19'b0000000_111011101101;
      15'b001_001001100011 : VALUE=19'b0000000_111011101101;
      15'b001_001001100100 : VALUE=19'b0000000_111011101101;
      15'b001_001001100101 : VALUE=19'b0000000_111011101100;
      15'b001_001001100110 : VALUE=19'b0000000_111011101100;
      15'b001_001001100111 : VALUE=19'b0000000_111011101011;
      15'b001_001001101000 : VALUE=19'b0000000_111011101011;
      15'b001_001001101001 : VALUE=19'b0000000_111011101010;
      15'b001_001001101010 : VALUE=19'b0000000_111011101010;
      15'b001_001001101011 : VALUE=19'b0000000_111011101010;
      15'b001_001001101100 : VALUE=19'b0000000_111011101001;
      15'b001_001001101101 : VALUE=19'b0000000_111011101001;
      15'b001_001001101110 : VALUE=19'b0000000_111011101000;
      15'b001_001001101111 : VALUE=19'b0000000_111011101000;
      15'b001_001001110000 : VALUE=19'b0000000_111011101000;
      15'b001_001001110001 : VALUE=19'b0000000_111011100111;
      15'b001_001001110010 : VALUE=19'b0000000_111011100111;
      15'b001_001001110011 : VALUE=19'b0000000_111011100110;
      15'b001_001001110100 : VALUE=19'b0000000_111011100110;
      15'b001_001001110101 : VALUE=19'b0000000_111011100110;
      15'b001_001001110110 : VALUE=19'b0000000_111011100101;
      15'b001_001001110111 : VALUE=19'b0000000_111011100101;
      15'b001_001001111000 : VALUE=19'b0000000_111011100100;
      15'b001_001001111001 : VALUE=19'b0000000_111011100100;
      15'b001_001001111010 : VALUE=19'b0000000_111011100100;
      15'b001_001001111011 : VALUE=19'b0000000_111011100011;
      15'b001_001001111100 : VALUE=19'b0000000_111011100011;
      15'b001_001001111101 : VALUE=19'b0000000_111011100010;
      15'b001_001001111110 : VALUE=19'b0000000_111011100010;
      15'b001_001001111111 : VALUE=19'b0000000_111011100010;
      15'b001_001010000000 : VALUE=19'b0000000_111011100001;
      15'b001_001010000001 : VALUE=19'b0000000_111011100001;
      15'b001_001010000010 : VALUE=19'b0000000_111011100000;
      15'b001_001010000011 : VALUE=19'b0000000_111011100000;
      15'b001_001010000100 : VALUE=19'b0000000_111011100000;
      15'b001_001010000101 : VALUE=19'b0000000_111011011111;
      15'b001_001010000110 : VALUE=19'b0000000_111011011111;
      15'b001_001010000111 : VALUE=19'b0000000_111011011110;
      15'b001_001010001000 : VALUE=19'b0000000_111011011110;
      15'b001_001010001001 : VALUE=19'b0000000_111011011110;
      15'b001_001010001010 : VALUE=19'b0000000_111011011101;
      15'b001_001010001011 : VALUE=19'b0000000_111011011101;
      15'b001_001010001100 : VALUE=19'b0000000_111011011100;
      15'b001_001010001101 : VALUE=19'b0000000_111011011100;
      15'b001_001010001110 : VALUE=19'b0000000_111011011100;
      15'b001_001010001111 : VALUE=19'b0000000_111011011011;
      15'b001_001010010000 : VALUE=19'b0000000_111011011011;
      15'b001_001010010001 : VALUE=19'b0000000_111011011010;
      15'b001_001010010010 : VALUE=19'b0000000_111011011010;
      15'b001_001010010011 : VALUE=19'b0000000_111011011010;
      15'b001_001010010100 : VALUE=19'b0000000_111011011001;
      15'b001_001010010101 : VALUE=19'b0000000_111011011001;
      15'b001_001010010110 : VALUE=19'b0000000_111011011000;
      15'b001_001010010111 : VALUE=19'b0000000_111011011000;
      15'b001_001010011000 : VALUE=19'b0000000_111011011000;
      15'b001_001010011001 : VALUE=19'b0000000_111011010111;
      15'b001_001010011010 : VALUE=19'b0000000_111011010111;
      15'b001_001010011011 : VALUE=19'b0000000_111011010110;
      15'b001_001010011100 : VALUE=19'b0000000_111011010110;
      15'b001_001010011101 : VALUE=19'b0000000_111011010110;
      15'b001_001010011110 : VALUE=19'b0000000_111011010101;
      15'b001_001010011111 : VALUE=19'b0000000_111011010101;
      15'b001_001010100000 : VALUE=19'b0000000_111011010100;
      15'b001_001010100001 : VALUE=19'b0000000_111011010100;
      15'b001_001010100010 : VALUE=19'b0000000_111011010100;
      15'b001_001010100011 : VALUE=19'b0000000_111011010011;
      15'b001_001010100100 : VALUE=19'b0000000_111011010011;
      15'b001_001010100101 : VALUE=19'b0000000_111011010010;
      15'b001_001010100110 : VALUE=19'b0000000_111011010010;
      15'b001_001010100111 : VALUE=19'b0000000_111011010010;
      15'b001_001010101000 : VALUE=19'b0000000_111011010001;
      15'b001_001010101001 : VALUE=19'b0000000_111011010001;
      15'b001_001010101010 : VALUE=19'b0000000_111011010000;
      15'b001_001010101011 : VALUE=19'b0000000_111011010000;
      15'b001_001010101100 : VALUE=19'b0000000_111011010000;
      15'b001_001010101101 : VALUE=19'b0000000_111011001111;
      15'b001_001010101110 : VALUE=19'b0000000_111011001111;
      15'b001_001010101111 : VALUE=19'b0000000_111011001110;
      15'b001_001010110000 : VALUE=19'b0000000_111011001110;
      15'b001_001010110001 : VALUE=19'b0000000_111011001110;
      15'b001_001010110010 : VALUE=19'b0000000_111011001101;
      15'b001_001010110011 : VALUE=19'b0000000_111011001101;
      15'b001_001010110100 : VALUE=19'b0000000_111011001100;
      15'b001_001010110101 : VALUE=19'b0000000_111011001100;
      15'b001_001010110110 : VALUE=19'b0000000_111011001100;
      15'b001_001010110111 : VALUE=19'b0000000_111011001011;
      15'b001_001010111000 : VALUE=19'b0000000_111011001011;
      15'b001_001010111001 : VALUE=19'b0000000_111011001010;
      15'b001_001010111010 : VALUE=19'b0000000_111011001010;
      15'b001_001010111011 : VALUE=19'b0000000_111011001010;
      15'b001_001010111100 : VALUE=19'b0000000_111011001001;
      15'b001_001010111101 : VALUE=19'b0000000_111011001001;
      15'b001_001010111110 : VALUE=19'b0000000_111011001001;
      15'b001_001010111111 : VALUE=19'b0000000_111011001000;
      15'b001_001011000000 : VALUE=19'b0000000_111011001000;
      15'b001_001011000001 : VALUE=19'b0000000_111011000111;
      15'b001_001011000010 : VALUE=19'b0000000_111011000111;
      15'b001_001011000011 : VALUE=19'b0000000_111011000111;
      15'b001_001011000100 : VALUE=19'b0000000_111011000110;
      15'b001_001011000101 : VALUE=19'b0000000_111011000110;
      15'b001_001011000110 : VALUE=19'b0000000_111011000101;
      15'b001_001011000111 : VALUE=19'b0000000_111011000101;
      15'b001_001011001000 : VALUE=19'b0000000_111011000101;
      15'b001_001011001001 : VALUE=19'b0000000_111011000100;
      15'b001_001011001010 : VALUE=19'b0000000_111011000100;
      15'b001_001011001011 : VALUE=19'b0000000_111011000011;
      15'b001_001011001100 : VALUE=19'b0000000_111011000011;
      15'b001_001011001101 : VALUE=19'b0000000_111011000011;
      15'b001_001011001110 : VALUE=19'b0000000_111011000010;
      15'b001_001011001111 : VALUE=19'b0000000_111011000010;
      15'b001_001011010000 : VALUE=19'b0000000_111011000001;
      15'b001_001011010001 : VALUE=19'b0000000_111011000001;
      15'b001_001011010010 : VALUE=19'b0000000_111011000001;
      15'b001_001011010011 : VALUE=19'b0000000_111011000000;
      15'b001_001011010100 : VALUE=19'b0000000_111011000000;
      15'b001_001011010101 : VALUE=19'b0000000_111010111111;
      15'b001_001011010110 : VALUE=19'b0000000_111010111111;
      15'b001_001011010111 : VALUE=19'b0000000_111010111111;
      15'b001_001011011000 : VALUE=19'b0000000_111010111110;
      15'b001_001011011001 : VALUE=19'b0000000_111010111110;
      15'b001_001011011010 : VALUE=19'b0000000_111010111110;
      15'b001_001011011011 : VALUE=19'b0000000_111010111101;
      15'b001_001011011100 : VALUE=19'b0000000_111010111101;
      15'b001_001011011101 : VALUE=19'b0000000_111010111100;
      15'b001_001011011110 : VALUE=19'b0000000_111010111100;
      15'b001_001011011111 : VALUE=19'b0000000_111010111100;
      15'b001_001011100000 : VALUE=19'b0000000_111010111011;
      15'b001_001011100001 : VALUE=19'b0000000_111010111011;
      15'b001_001011100010 : VALUE=19'b0000000_111010111010;
      15'b001_001011100011 : VALUE=19'b0000000_111010111010;
      15'b001_001011100100 : VALUE=19'b0000000_111010111010;
      15'b001_001011100101 : VALUE=19'b0000000_111010111001;
      15'b001_001011100110 : VALUE=19'b0000000_111010111001;
      15'b001_001011100111 : VALUE=19'b0000000_111010111000;
      15'b001_001011101000 : VALUE=19'b0000000_111010111000;
      15'b001_001011101001 : VALUE=19'b0000000_111010111000;
      15'b001_001011101010 : VALUE=19'b0000000_111010110111;
      15'b001_001011101011 : VALUE=19'b0000000_111010110111;
      15'b001_001011101100 : VALUE=19'b0000000_111010110110;
      15'b001_001011101101 : VALUE=19'b0000000_111010110110;
      15'b001_001011101110 : VALUE=19'b0000000_111010110110;
      15'b001_001011101111 : VALUE=19'b0000000_111010110101;
      15'b001_001011110000 : VALUE=19'b0000000_111010110101;
      15'b001_001011110001 : VALUE=19'b0000000_111010110101;
      15'b001_001011110010 : VALUE=19'b0000000_111010110100;
      15'b001_001011110011 : VALUE=19'b0000000_111010110100;
      15'b001_001011110100 : VALUE=19'b0000000_111010110011;
      15'b001_001011110101 : VALUE=19'b0000000_111010110011;
      15'b001_001011110110 : VALUE=19'b0000000_111010110011;
      15'b001_001011110111 : VALUE=19'b0000000_111010110010;
      15'b001_001011111000 : VALUE=19'b0000000_111010110010;
      15'b001_001011111001 : VALUE=19'b0000000_111010110001;
      15'b001_001011111010 : VALUE=19'b0000000_111010110001;
      15'b001_001011111011 : VALUE=19'b0000000_111010110001;
      15'b001_001011111100 : VALUE=19'b0000000_111010110000;
      15'b001_001011111101 : VALUE=19'b0000000_111010110000;
      15'b001_001011111110 : VALUE=19'b0000000_111010110000;
      15'b001_001011111111 : VALUE=19'b0000000_111010101111;
      15'b001_001100000000 : VALUE=19'b0000000_111010101111;
      15'b001_001100000001 : VALUE=19'b0000000_111010101110;
      15'b001_001100000010 : VALUE=19'b0000000_111010101110;
      15'b001_001100000011 : VALUE=19'b0000000_111010101110;
      15'b001_001100000100 : VALUE=19'b0000000_111010101101;
      15'b001_001100000101 : VALUE=19'b0000000_111010101101;
      15'b001_001100000110 : VALUE=19'b0000000_111010101100;
      15'b001_001100000111 : VALUE=19'b0000000_111010101100;
      15'b001_001100001000 : VALUE=19'b0000000_111010101100;
      15'b001_001100001001 : VALUE=19'b0000000_111010101011;
      15'b001_001100001010 : VALUE=19'b0000000_111010101011;
      15'b001_001100001011 : VALUE=19'b0000000_111010101011;
      15'b001_001100001100 : VALUE=19'b0000000_111010101010;
      15'b001_001100001101 : VALUE=19'b0000000_111010101010;
      15'b001_001100001110 : VALUE=19'b0000000_111010101001;
      15'b001_001100001111 : VALUE=19'b0000000_111010101001;
      15'b001_001100010000 : VALUE=19'b0000000_111010101001;
      15'b001_001100010001 : VALUE=19'b0000000_111010101000;
      15'b001_001100010010 : VALUE=19'b0000000_111010101000;
      15'b001_001100010011 : VALUE=19'b0000000_111010100111;
      15'b001_001100010100 : VALUE=19'b0000000_111010100111;
      15'b001_001100010101 : VALUE=19'b0000000_111010100111;
      15'b001_001100010110 : VALUE=19'b0000000_111010100110;
      15'b001_001100010111 : VALUE=19'b0000000_111010100110;
      15'b001_001100011000 : VALUE=19'b0000000_111010100110;
      15'b001_001100011001 : VALUE=19'b0000000_111010100101;
      15'b001_001100011010 : VALUE=19'b0000000_111010100101;
      15'b001_001100011011 : VALUE=19'b0000000_111010100100;
      15'b001_001100011100 : VALUE=19'b0000000_111010100100;
      15'b001_001100011101 : VALUE=19'b0000000_111010100100;
      15'b001_001100011110 : VALUE=19'b0000000_111010100011;
      15'b001_001100011111 : VALUE=19'b0000000_111010100011;
      15'b001_001100100000 : VALUE=19'b0000000_111010100010;
      15'b001_001100100001 : VALUE=19'b0000000_111010100010;
      15'b001_001100100010 : VALUE=19'b0000000_111010100010;
      15'b001_001100100011 : VALUE=19'b0000000_111010100001;
      15'b001_001100100100 : VALUE=19'b0000000_111010100001;
      15'b001_001100100101 : VALUE=19'b0000000_111010100001;
      15'b001_001100100110 : VALUE=19'b0000000_111010100000;
      15'b001_001100100111 : VALUE=19'b0000000_111010100000;
      15'b001_001100101000 : VALUE=19'b0000000_111010011111;
      15'b001_001100101001 : VALUE=19'b0000000_111010011111;
      15'b001_001100101010 : VALUE=19'b0000000_111010011111;
      15'b001_001100101011 : VALUE=19'b0000000_111010011110;
      15'b001_001100101100 : VALUE=19'b0000000_111010011110;
      15'b001_001100101101 : VALUE=19'b0000000_111010011101;
      15'b001_001100101110 : VALUE=19'b0000000_111010011101;
      15'b001_001100101111 : VALUE=19'b0000000_111010011101;
      15'b001_001100110000 : VALUE=19'b0000000_111010011100;
      15'b001_001100110001 : VALUE=19'b0000000_111010011100;
      15'b001_001100110010 : VALUE=19'b0000000_111010011100;
      15'b001_001100110011 : VALUE=19'b0000000_111010011011;
      15'b001_001100110100 : VALUE=19'b0000000_111010011011;
      15'b001_001100110101 : VALUE=19'b0000000_111010011010;
      15'b001_001100110110 : VALUE=19'b0000000_111010011010;
      15'b001_001100110111 : VALUE=19'b0000000_111010011010;
      15'b001_001100111000 : VALUE=19'b0000000_111010011001;
      15'b001_001100111001 : VALUE=19'b0000000_111010011001;
      15'b001_001100111010 : VALUE=19'b0000000_111010011001;
      15'b001_001100111011 : VALUE=19'b0000000_111010011000;
      15'b001_001100111100 : VALUE=19'b0000000_111010011000;
      15'b001_001100111101 : VALUE=19'b0000000_111010010111;
      15'b001_001100111110 : VALUE=19'b0000000_111010010111;
      15'b001_001100111111 : VALUE=19'b0000000_111010010111;
      15'b001_001101000000 : VALUE=19'b0000000_111010010110;
      15'b001_001101000001 : VALUE=19'b0000000_111010010110;
      15'b001_001101000010 : VALUE=19'b0000000_111010010110;
      15'b001_001101000011 : VALUE=19'b0000000_111010010101;
      15'b001_001101000100 : VALUE=19'b0000000_111010010101;
      15'b001_001101000101 : VALUE=19'b0000000_111010010100;
      15'b001_001101000110 : VALUE=19'b0000000_111010010100;
      15'b001_001101000111 : VALUE=19'b0000000_111010010100;
      15'b001_001101001000 : VALUE=19'b0000000_111010010011;
      15'b001_001101001001 : VALUE=19'b0000000_111010010011;
      15'b001_001101001010 : VALUE=19'b0000000_111010010010;
      15'b001_001101001011 : VALUE=19'b0000000_111010010010;
      15'b001_001101001100 : VALUE=19'b0000000_111010010010;
      15'b001_001101001101 : VALUE=19'b0000000_111010010001;
      15'b001_001101001110 : VALUE=19'b0000000_111010010001;
      15'b001_001101001111 : VALUE=19'b0000000_111010010001;
      15'b001_001101010000 : VALUE=19'b0000000_111010010000;
      15'b001_001101010001 : VALUE=19'b0000000_111010010000;
      15'b001_001101010010 : VALUE=19'b0000000_111010001111;
      15'b001_001101010011 : VALUE=19'b0000000_111010001111;
      15'b001_001101010100 : VALUE=19'b0000000_111010001111;
      15'b001_001101010101 : VALUE=19'b0000000_111010001110;
      15'b001_001101010110 : VALUE=19'b0000000_111010001110;
      15'b001_001101010111 : VALUE=19'b0000000_111010001110;
      15'b001_001101011000 : VALUE=19'b0000000_111010001101;
      15'b001_001101011001 : VALUE=19'b0000000_111010001101;
      15'b001_001101011010 : VALUE=19'b0000000_111010001100;
      15'b001_001101011011 : VALUE=19'b0000000_111010001100;
      15'b001_001101011100 : VALUE=19'b0000000_111010001100;
      15'b001_001101011101 : VALUE=19'b0000000_111010001011;
      15'b001_001101011110 : VALUE=19'b0000000_111010001011;
      15'b001_001101011111 : VALUE=19'b0000000_111010001011;
      15'b001_001101100000 : VALUE=19'b0000000_111010001010;
      15'b001_001101100001 : VALUE=19'b0000000_111010001010;
      15'b001_001101100010 : VALUE=19'b0000000_111010001001;
      15'b001_001101100011 : VALUE=19'b0000000_111010001001;
      15'b001_001101100100 : VALUE=19'b0000000_111010001001;
      15'b001_001101100101 : VALUE=19'b0000000_111010001000;
      15'b001_001101100110 : VALUE=19'b0000000_111010001000;
      15'b001_001101100111 : VALUE=19'b0000000_111010001000;
      15'b001_001101101000 : VALUE=19'b0000000_111010000111;
      15'b001_001101101001 : VALUE=19'b0000000_111010000111;
      15'b001_001101101010 : VALUE=19'b0000000_111010000110;
      15'b001_001101101011 : VALUE=19'b0000000_111010000110;
      15'b001_001101101100 : VALUE=19'b0000000_111010000110;
      15'b001_001101101101 : VALUE=19'b0000000_111010000101;
      15'b001_001101101110 : VALUE=19'b0000000_111010000101;
      15'b001_001101101111 : VALUE=19'b0000000_111010000101;
      15'b001_001101110000 : VALUE=19'b0000000_111010000100;
      15'b001_001101110001 : VALUE=19'b0000000_111010000100;
      15'b001_001101110010 : VALUE=19'b0000000_111010000011;
      15'b001_001101110011 : VALUE=19'b0000000_111010000011;
      15'b001_001101110100 : VALUE=19'b0000000_111010000011;
      15'b001_001101110101 : VALUE=19'b0000000_111010000010;
      15'b001_001101110110 : VALUE=19'b0000000_111010000010;
      15'b001_001101110111 : VALUE=19'b0000000_111010000010;
      15'b001_001101111000 : VALUE=19'b0000000_111010000001;
      15'b001_001101111001 : VALUE=19'b0000000_111010000001;
      15'b001_001101111010 : VALUE=19'b0000000_111010000000;
      15'b001_001101111011 : VALUE=19'b0000000_111010000000;
      15'b001_001101111100 : VALUE=19'b0000000_111010000000;
      15'b001_001101111101 : VALUE=19'b0000000_111001111111;
      15'b001_001101111110 : VALUE=19'b0000000_111001111111;
      15'b001_001101111111 : VALUE=19'b0000000_111001111111;
      15'b001_001110000000 : VALUE=19'b0000000_111001111110;
      15'b001_001110000001 : VALUE=19'b0000000_111001111110;
      15'b001_001110000010 : VALUE=19'b0000000_111001111110;
      15'b001_001110000011 : VALUE=19'b0000000_111001111101;
      15'b001_001110000100 : VALUE=19'b0000000_111001111101;
      15'b001_001110000101 : VALUE=19'b0000000_111001111100;
      15'b001_001110000110 : VALUE=19'b0000000_111001111100;
      15'b001_001110000111 : VALUE=19'b0000000_111001111100;
      15'b001_001110001000 : VALUE=19'b0000000_111001111011;
      15'b001_001110001001 : VALUE=19'b0000000_111001111011;
      15'b001_001110001010 : VALUE=19'b0000000_111001111011;
      15'b001_001110001011 : VALUE=19'b0000000_111001111010;
      15'b001_001110001100 : VALUE=19'b0000000_111001111010;
      15'b001_001110001101 : VALUE=19'b0000000_111001111001;
      15'b001_001110001110 : VALUE=19'b0000000_111001111001;
      15'b001_001110001111 : VALUE=19'b0000000_111001111001;
      15'b001_001110010000 : VALUE=19'b0000000_111001111000;
      15'b001_001110010001 : VALUE=19'b0000000_111001111000;
      15'b001_001110010010 : VALUE=19'b0000000_111001111000;
      15'b001_001110010011 : VALUE=19'b0000000_111001110111;
      15'b001_001110010100 : VALUE=19'b0000000_111001110111;
      15'b001_001110010101 : VALUE=19'b0000000_111001110110;
      15'b001_001110010110 : VALUE=19'b0000000_111001110110;
      15'b001_001110010111 : VALUE=19'b0000000_111001110110;
      15'b001_001110011000 : VALUE=19'b0000000_111001110101;
      15'b001_001110011001 : VALUE=19'b0000000_111001110101;
      15'b001_001110011010 : VALUE=19'b0000000_111001110101;
      15'b001_001110011011 : VALUE=19'b0000000_111001110100;
      15'b001_001110011100 : VALUE=19'b0000000_111001110100;
      15'b001_001110011101 : VALUE=19'b0000000_111001110100;
      15'b001_001110011110 : VALUE=19'b0000000_111001110011;
      15'b001_001110011111 : VALUE=19'b0000000_111001110011;
      15'b001_001110100000 : VALUE=19'b0000000_111001110010;
      15'b001_001110100001 : VALUE=19'b0000000_111001110010;
      15'b001_001110100010 : VALUE=19'b0000000_111001110010;
      15'b001_001110100011 : VALUE=19'b0000000_111001110001;
      15'b001_001110100100 : VALUE=19'b0000000_111001110001;
      15'b001_001110100101 : VALUE=19'b0000000_111001110001;
      15'b001_001110100110 : VALUE=19'b0000000_111001110000;
      15'b001_001110100111 : VALUE=19'b0000000_111001110000;
      15'b001_001110101000 : VALUE=19'b0000000_111001101111;
      15'b001_001110101001 : VALUE=19'b0000000_111001101111;
      15'b001_001110101010 : VALUE=19'b0000000_111001101111;
      15'b001_001110101011 : VALUE=19'b0000000_111001101110;
      15'b001_001110101100 : VALUE=19'b0000000_111001101110;
      15'b001_001110101101 : VALUE=19'b0000000_111001101110;
      15'b001_001110101110 : VALUE=19'b0000000_111001101101;
      15'b001_001110101111 : VALUE=19'b0000000_111001101101;
      15'b001_001110110000 : VALUE=19'b0000000_111001101101;
      15'b001_001110110001 : VALUE=19'b0000000_111001101100;
      15'b001_001110110010 : VALUE=19'b0000000_111001101100;
      15'b001_001110110011 : VALUE=19'b0000000_111001101011;
      15'b001_001110110100 : VALUE=19'b0000000_111001101011;
      15'b001_001110110101 : VALUE=19'b0000000_111001101011;
      15'b001_001110110110 : VALUE=19'b0000000_111001101010;
      15'b001_001110110111 : VALUE=19'b0000000_111001101010;
      15'b001_001110111000 : VALUE=19'b0000000_111001101010;
      15'b001_001110111001 : VALUE=19'b0000000_111001101001;
      15'b001_001110111010 : VALUE=19'b0000000_111001101001;
      15'b001_001110111011 : VALUE=19'b0000000_111001101001;
      15'b001_001110111100 : VALUE=19'b0000000_111001101000;
      15'b001_001110111101 : VALUE=19'b0000000_111001101000;
      15'b001_001110111110 : VALUE=19'b0000000_111001100111;
      15'b001_001110111111 : VALUE=19'b0000000_111001100111;
      15'b001_001111000000 : VALUE=19'b0000000_111001100111;
      15'b001_001111000001 : VALUE=19'b0000000_111001100110;
      15'b001_001111000010 : VALUE=19'b0000000_111001100110;
      15'b001_001111000011 : VALUE=19'b0000000_111001100110;
      15'b001_001111000100 : VALUE=19'b0000000_111001100101;
      15'b001_001111000101 : VALUE=19'b0000000_111001100101;
      15'b001_001111000110 : VALUE=19'b0000000_111001100101;
      15'b001_001111000111 : VALUE=19'b0000000_111001100100;
      15'b001_001111001000 : VALUE=19'b0000000_111001100100;
      15'b001_001111001001 : VALUE=19'b0000000_111001100011;
      15'b001_001111001010 : VALUE=19'b0000000_111001100011;
      15'b001_001111001011 : VALUE=19'b0000000_111001100011;
      15'b001_001111001100 : VALUE=19'b0000000_111001100010;
      15'b001_001111001101 : VALUE=19'b0000000_111001100010;
      15'b001_001111001110 : VALUE=19'b0000000_111001100010;
      15'b001_001111001111 : VALUE=19'b0000000_111001100001;
      15'b001_001111010000 : VALUE=19'b0000000_111001100001;
      15'b001_001111010001 : VALUE=19'b0000000_111001100001;
      15'b001_001111010010 : VALUE=19'b0000000_111001100000;
      15'b001_001111010011 : VALUE=19'b0000000_111001100000;
      15'b001_001111010100 : VALUE=19'b0000000_111001011111;
      15'b001_001111010101 : VALUE=19'b0000000_111001011111;
      15'b001_001111010110 : VALUE=19'b0000000_111001011111;
      15'b001_001111010111 : VALUE=19'b0000000_111001011110;
      15'b001_001111011000 : VALUE=19'b0000000_111001011110;
      15'b001_001111011001 : VALUE=19'b0000000_111001011110;
      15'b001_001111011010 : VALUE=19'b0000000_111001011101;
      15'b001_001111011011 : VALUE=19'b0000000_111001011101;
      15'b001_001111011100 : VALUE=19'b0000000_111001011101;
      15'b001_001111011101 : VALUE=19'b0000000_111001011100;
      15'b001_001111011110 : VALUE=19'b0000000_111001011100;
      15'b001_001111011111 : VALUE=19'b0000000_111001011011;
      15'b001_001111100000 : VALUE=19'b0000000_111001011011;
      15'b001_001111100001 : VALUE=19'b0000000_111001011011;
      15'b001_001111100010 : VALUE=19'b0000000_111001011010;
      15'b001_001111100011 : VALUE=19'b0000000_111001011010;
      15'b001_001111100100 : VALUE=19'b0000000_111001011010;
      15'b001_001111100101 : VALUE=19'b0000000_111001011001;
      15'b001_001111100110 : VALUE=19'b0000000_111001011001;
      15'b001_001111100111 : VALUE=19'b0000000_111001011001;
      15'b001_001111101000 : VALUE=19'b0000000_111001011000;
      15'b001_001111101001 : VALUE=19'b0000000_111001011000;
      15'b001_001111101010 : VALUE=19'b0000000_111001010111;
      15'b001_001111101011 : VALUE=19'b0000000_111001010111;
      15'b001_001111101100 : VALUE=19'b0000000_111001010111;
      15'b001_001111101101 : VALUE=19'b0000000_111001010110;
      15'b001_001111101110 : VALUE=19'b0000000_111001010110;
      15'b001_001111101111 : VALUE=19'b0000000_111001010110;
      15'b001_001111110000 : VALUE=19'b0000000_111001010101;
      15'b001_001111110001 : VALUE=19'b0000000_111001010101;
      15'b001_001111110010 : VALUE=19'b0000000_111001010101;
      15'b001_001111110011 : VALUE=19'b0000000_111001010100;
      15'b001_001111110100 : VALUE=19'b0000000_111001010100;
      15'b001_001111110101 : VALUE=19'b0000000_111001010100;
      15'b001_001111110110 : VALUE=19'b0000000_111001010011;
      15'b001_001111110111 : VALUE=19'b0000000_111001010011;
      15'b001_001111111000 : VALUE=19'b0000000_111001010010;
      15'b001_001111111001 : VALUE=19'b0000000_111001010010;
      15'b001_001111111010 : VALUE=19'b0000000_111001010010;
      15'b001_001111111011 : VALUE=19'b0000000_111001010001;
      15'b001_001111111100 : VALUE=19'b0000000_111001010001;
      15'b001_001111111101 : VALUE=19'b0000000_111001010001;
      15'b001_001111111110 : VALUE=19'b0000000_111001010000;
      15'b001_001111111111 : VALUE=19'b0000000_111001010000;
      15'b001_010000000000 : VALUE=19'b0000000_111001010000;
      15'b001_010000000001 : VALUE=19'b0000000_111001001111;
      15'b001_010000000010 : VALUE=19'b0000000_111001001111;
      15'b001_010000000011 : VALUE=19'b0000000_111001001111;
      15'b001_010000000100 : VALUE=19'b0000000_111001001110;
      15'b001_010000000101 : VALUE=19'b0000000_111001001110;
      15'b001_010000000110 : VALUE=19'b0000000_111001001101;
      15'b001_010000000111 : VALUE=19'b0000000_111001001101;
      15'b001_010000001000 : VALUE=19'b0000000_111001001101;
      15'b001_010000001001 : VALUE=19'b0000000_111001001100;
      15'b001_010000001010 : VALUE=19'b0000000_111001001100;
      15'b001_010000001011 : VALUE=19'b0000000_111001001100;
      15'b001_010000001100 : VALUE=19'b0000000_111001001011;
      15'b001_010000001101 : VALUE=19'b0000000_111001001011;
      15'b001_010000001110 : VALUE=19'b0000000_111001001011;
      15'b001_010000001111 : VALUE=19'b0000000_111001001010;
      15'b001_010000010000 : VALUE=19'b0000000_111001001010;
      15'b001_010000010001 : VALUE=19'b0000000_111001001010;
      15'b001_010000010010 : VALUE=19'b0000000_111001001001;
      15'b001_010000010011 : VALUE=19'b0000000_111001001001;
      15'b001_010000010100 : VALUE=19'b0000000_111001001000;
      15'b001_010000010101 : VALUE=19'b0000000_111001001000;
      15'b001_010000010110 : VALUE=19'b0000000_111001001000;
      15'b001_010000010111 : VALUE=19'b0000000_111001000111;
      15'b001_010000011000 : VALUE=19'b0000000_111001000111;
      15'b001_010000011001 : VALUE=19'b0000000_111001000111;
      15'b001_010000011010 : VALUE=19'b0000000_111001000110;
      15'b001_010000011011 : VALUE=19'b0000000_111001000110;
      15'b001_010000011100 : VALUE=19'b0000000_111001000110;
      15'b001_010000011101 : VALUE=19'b0000000_111001000101;
      15'b001_010000011110 : VALUE=19'b0000000_111001000101;
      15'b001_010000011111 : VALUE=19'b0000000_111001000101;
      15'b001_010000100000 : VALUE=19'b0000000_111001000100;
      15'b001_010000100001 : VALUE=19'b0000000_111001000100;
      15'b001_010000100010 : VALUE=19'b0000000_111001000011;
      15'b001_010000100011 : VALUE=19'b0000000_111001000011;
      15'b001_010000100100 : VALUE=19'b0000000_111001000011;
      15'b001_010000100101 : VALUE=19'b0000000_111001000010;
      15'b001_010000100110 : VALUE=19'b0000000_111001000010;
      15'b001_010000100111 : VALUE=19'b0000000_111001000010;
      15'b001_010000101000 : VALUE=19'b0000000_111001000001;
      15'b001_010000101001 : VALUE=19'b0000000_111001000001;
      15'b001_010000101010 : VALUE=19'b0000000_111001000001;
      15'b001_010000101011 : VALUE=19'b0000000_111001000000;
      15'b001_010000101100 : VALUE=19'b0000000_111001000000;
      15'b001_010000101101 : VALUE=19'b0000000_111001000000;
      15'b001_010000101110 : VALUE=19'b0000000_111000111111;
      15'b001_010000101111 : VALUE=19'b0000000_111000111111;
      15'b001_010000110000 : VALUE=19'b0000000_111000111111;
      15'b001_010000110001 : VALUE=19'b0000000_111000111110;
      15'b001_010000110010 : VALUE=19'b0000000_111000111110;
      15'b001_010000110011 : VALUE=19'b0000000_111000111101;
      15'b001_010000110100 : VALUE=19'b0000000_111000111101;
      15'b001_010000110101 : VALUE=19'b0000000_111000111101;
      15'b001_010000110110 : VALUE=19'b0000000_111000111100;
      15'b001_010000110111 : VALUE=19'b0000000_111000111100;
      15'b001_010000111000 : VALUE=19'b0000000_111000111100;
      15'b001_010000111001 : VALUE=19'b0000000_111000111011;
      15'b001_010000111010 : VALUE=19'b0000000_111000111011;
      15'b001_010000111011 : VALUE=19'b0000000_111000111011;
      15'b001_010000111100 : VALUE=19'b0000000_111000111010;
      15'b001_010000111101 : VALUE=19'b0000000_111000111010;
      15'b001_010000111110 : VALUE=19'b0000000_111000111010;
      15'b001_010000111111 : VALUE=19'b0000000_111000111001;
      15'b001_010001000000 : VALUE=19'b0000000_111000111001;
      15'b001_010001000001 : VALUE=19'b0000000_111000111001;
      15'b001_010001000010 : VALUE=19'b0000000_111000111000;
      15'b001_010001000011 : VALUE=19'b0000000_111000111000;
      15'b001_010001000100 : VALUE=19'b0000000_111000110111;
      15'b001_010001000101 : VALUE=19'b0000000_111000110111;
      15'b001_010001000110 : VALUE=19'b0000000_111000110111;
      15'b001_010001000111 : VALUE=19'b0000000_111000110110;
      15'b001_010001001000 : VALUE=19'b0000000_111000110110;
      15'b001_010001001001 : VALUE=19'b0000000_111000110110;
      15'b001_010001001010 : VALUE=19'b0000000_111000110101;
      15'b001_010001001011 : VALUE=19'b0000000_111000110101;
      15'b001_010001001100 : VALUE=19'b0000000_111000110101;
      15'b001_010001001101 : VALUE=19'b0000000_111000110100;
      15'b001_010001001110 : VALUE=19'b0000000_111000110100;
      15'b001_010001001111 : VALUE=19'b0000000_111000110100;
      15'b001_010001010000 : VALUE=19'b0000000_111000110011;
      15'b001_010001010001 : VALUE=19'b0000000_111000110011;
      15'b001_010001010010 : VALUE=19'b0000000_111000110011;
      15'b001_010001010011 : VALUE=19'b0000000_111000110010;
      15'b001_010001010100 : VALUE=19'b0000000_111000110010;
      15'b001_010001010101 : VALUE=19'b0000000_111000110010;
      15'b001_010001010110 : VALUE=19'b0000000_111000110001;
      15'b001_010001010111 : VALUE=19'b0000000_111000110001;
      15'b001_010001011000 : VALUE=19'b0000000_111000110000;
      15'b001_010001011001 : VALUE=19'b0000000_111000110000;
      15'b001_010001011010 : VALUE=19'b0000000_111000110000;
      15'b001_010001011011 : VALUE=19'b0000000_111000101111;
      15'b001_010001011100 : VALUE=19'b0000000_111000101111;
      15'b001_010001011101 : VALUE=19'b0000000_111000101111;
      15'b001_010001011110 : VALUE=19'b0000000_111000101110;
      15'b001_010001011111 : VALUE=19'b0000000_111000101110;
      15'b001_010001100000 : VALUE=19'b0000000_111000101110;
      15'b001_010001100001 : VALUE=19'b0000000_111000101101;
      15'b001_010001100010 : VALUE=19'b0000000_111000101101;
      15'b001_010001100011 : VALUE=19'b0000000_111000101101;
      15'b001_010001100100 : VALUE=19'b0000000_111000101100;
      15'b001_010001100101 : VALUE=19'b0000000_111000101100;
      15'b001_010001100110 : VALUE=19'b0000000_111000101100;
      15'b001_010001100111 : VALUE=19'b0000000_111000101011;
      15'b001_010001101000 : VALUE=19'b0000000_111000101011;
      15'b001_010001101001 : VALUE=19'b0000000_111000101011;
      15'b001_010001101010 : VALUE=19'b0000000_111000101010;
      15'b001_010001101011 : VALUE=19'b0000000_111000101010;
      15'b001_010001101100 : VALUE=19'b0000000_111000101010;
      15'b001_010001101101 : VALUE=19'b0000000_111000101001;
      15'b001_010001101110 : VALUE=19'b0000000_111000101001;
      15'b001_010001101111 : VALUE=19'b0000000_111000101000;
      15'b001_010001110000 : VALUE=19'b0000000_111000101000;
      15'b001_010001110001 : VALUE=19'b0000000_111000101000;
      15'b001_010001110010 : VALUE=19'b0000000_111000100111;
      15'b001_010001110011 : VALUE=19'b0000000_111000100111;
      15'b001_010001110100 : VALUE=19'b0000000_111000100111;
      15'b001_010001110101 : VALUE=19'b0000000_111000100110;
      15'b001_010001110110 : VALUE=19'b0000000_111000100110;
      15'b001_010001110111 : VALUE=19'b0000000_111000100110;
      15'b001_010001111000 : VALUE=19'b0000000_111000100101;
      15'b001_010001111001 : VALUE=19'b0000000_111000100101;
      15'b001_010001111010 : VALUE=19'b0000000_111000100101;
      15'b001_010001111011 : VALUE=19'b0000000_111000100100;
      15'b001_010001111100 : VALUE=19'b0000000_111000100100;
      15'b001_010001111101 : VALUE=19'b0000000_111000100100;
      15'b001_010001111110 : VALUE=19'b0000000_111000100011;
      15'b001_010001111111 : VALUE=19'b0000000_111000100011;
      15'b001_010010000000 : VALUE=19'b0000000_111000100011;
      15'b001_010010000001 : VALUE=19'b0000000_111000100010;
      15'b001_010010000010 : VALUE=19'b0000000_111000100010;
      15'b001_010010000011 : VALUE=19'b0000000_111000100010;
      15'b001_010010000100 : VALUE=19'b0000000_111000100001;
      15'b001_010010000101 : VALUE=19'b0000000_111000100001;
      15'b001_010010000110 : VALUE=19'b0000000_111000100001;
      15'b001_010010000111 : VALUE=19'b0000000_111000100000;
      15'b001_010010001000 : VALUE=19'b0000000_111000100000;
      15'b001_010010001001 : VALUE=19'b0000000_111000100000;
      15'b001_010010001010 : VALUE=19'b0000000_111000011111;
      15'b001_010010001011 : VALUE=19'b0000000_111000011111;
      15'b001_010010001100 : VALUE=19'b0000000_111000011110;
      15'b001_010010001101 : VALUE=19'b0000000_111000011110;
      15'b001_010010001110 : VALUE=19'b0000000_111000011110;
      15'b001_010010001111 : VALUE=19'b0000000_111000011101;
      15'b001_010010010000 : VALUE=19'b0000000_111000011101;
      15'b001_010010010001 : VALUE=19'b0000000_111000011101;
      15'b001_010010010010 : VALUE=19'b0000000_111000011100;
      15'b001_010010010011 : VALUE=19'b0000000_111000011100;
      15'b001_010010010100 : VALUE=19'b0000000_111000011100;
      15'b001_010010010101 : VALUE=19'b0000000_111000011011;
      15'b001_010010010110 : VALUE=19'b0000000_111000011011;
      15'b001_010010010111 : VALUE=19'b0000000_111000011011;
      15'b001_010010011000 : VALUE=19'b0000000_111000011010;
      15'b001_010010011001 : VALUE=19'b0000000_111000011010;
      15'b001_010010011010 : VALUE=19'b0000000_111000011010;
      15'b001_010010011011 : VALUE=19'b0000000_111000011001;
      15'b001_010010011100 : VALUE=19'b0000000_111000011001;
      15'b001_010010011101 : VALUE=19'b0000000_111000011001;
      15'b001_010010011110 : VALUE=19'b0000000_111000011000;
      15'b001_010010011111 : VALUE=19'b0000000_111000011000;
      15'b001_010010100000 : VALUE=19'b0000000_111000011000;
      15'b001_010010100001 : VALUE=19'b0000000_111000010111;
      15'b001_010010100010 : VALUE=19'b0000000_111000010111;
      15'b001_010010100011 : VALUE=19'b0000000_111000010111;
      15'b001_010010100100 : VALUE=19'b0000000_111000010110;
      15'b001_010010100101 : VALUE=19'b0000000_111000010110;
      15'b001_010010100110 : VALUE=19'b0000000_111000010110;
      15'b001_010010100111 : VALUE=19'b0000000_111000010101;
      15'b001_010010101000 : VALUE=19'b0000000_111000010101;
      15'b001_010010101001 : VALUE=19'b0000000_111000010101;
      15'b001_010010101010 : VALUE=19'b0000000_111000010100;
      15'b001_010010101011 : VALUE=19'b0000000_111000010100;
      15'b001_010010101100 : VALUE=19'b0000000_111000010100;
      15'b001_010010101101 : VALUE=19'b0000000_111000010011;
      15'b001_010010101110 : VALUE=19'b0000000_111000010011;
      15'b001_010010101111 : VALUE=19'b0000000_111000010011;
      15'b001_010010110000 : VALUE=19'b0000000_111000010010;
      15'b001_010010110001 : VALUE=19'b0000000_111000010010;
      15'b001_010010110010 : VALUE=19'b0000000_111000010010;
      15'b001_010010110011 : VALUE=19'b0000000_111000010001;
      15'b001_010010110100 : VALUE=19'b0000000_111000010001;
      15'b001_010010110101 : VALUE=19'b0000000_111000010000;
      15'b001_010010110110 : VALUE=19'b0000000_111000010000;
      15'b001_010010110111 : VALUE=19'b0000000_111000010000;
      15'b001_010010111000 : VALUE=19'b0000000_111000001111;
      15'b001_010010111001 : VALUE=19'b0000000_111000001111;
      15'b001_010010111010 : VALUE=19'b0000000_111000001111;
      15'b001_010010111011 : VALUE=19'b0000000_111000001110;
      15'b001_010010111100 : VALUE=19'b0000000_111000001110;
      15'b001_010010111101 : VALUE=19'b0000000_111000001110;
      15'b001_010010111110 : VALUE=19'b0000000_111000001101;
      15'b001_010010111111 : VALUE=19'b0000000_111000001101;
      15'b001_010011000000 : VALUE=19'b0000000_111000001101;
      15'b001_010011000001 : VALUE=19'b0000000_111000001100;
      15'b001_010011000010 : VALUE=19'b0000000_111000001100;
      15'b001_010011000011 : VALUE=19'b0000000_111000001100;
      15'b001_010011000100 : VALUE=19'b0000000_111000001011;
      15'b001_010011000101 : VALUE=19'b0000000_111000001011;
      15'b001_010011000110 : VALUE=19'b0000000_111000001011;
      15'b001_010011000111 : VALUE=19'b0000000_111000001010;
      15'b001_010011001000 : VALUE=19'b0000000_111000001010;
      15'b001_010011001001 : VALUE=19'b0000000_111000001010;
      15'b001_010011001010 : VALUE=19'b0000000_111000001001;
      15'b001_010011001011 : VALUE=19'b0000000_111000001001;
      15'b001_010011001100 : VALUE=19'b0000000_111000001001;
      15'b001_010011001101 : VALUE=19'b0000000_111000001000;
      15'b001_010011001110 : VALUE=19'b0000000_111000001000;
      15'b001_010011001111 : VALUE=19'b0000000_111000001000;
      15'b001_010011010000 : VALUE=19'b0000000_111000000111;
      15'b001_010011010001 : VALUE=19'b0000000_111000000111;
      15'b001_010011010010 : VALUE=19'b0000000_111000000111;
      15'b001_010011010011 : VALUE=19'b0000000_111000000110;
      15'b001_010011010100 : VALUE=19'b0000000_111000000110;
      15'b001_010011010101 : VALUE=19'b0000000_111000000110;
      15'b001_010011010110 : VALUE=19'b0000000_111000000101;
      15'b001_010011010111 : VALUE=19'b0000000_111000000101;
      15'b001_010011011000 : VALUE=19'b0000000_111000000101;
      15'b001_010011011001 : VALUE=19'b0000000_111000000100;
      15'b001_010011011010 : VALUE=19'b0000000_111000000100;
      15'b001_010011011011 : VALUE=19'b0000000_111000000100;
      15'b001_010011011100 : VALUE=19'b0000000_111000000011;
      15'b001_010011011101 : VALUE=19'b0000000_111000000011;
      15'b001_010011011110 : VALUE=19'b0000000_111000000011;
      15'b001_010011011111 : VALUE=19'b0000000_111000000010;
      15'b001_010011100000 : VALUE=19'b0000000_111000000010;
      15'b001_010011100001 : VALUE=19'b0000000_111000000010;
      15'b001_010011100010 : VALUE=19'b0000000_111000000001;
      15'b001_010011100011 : VALUE=19'b0000000_111000000001;
      15'b001_010011100100 : VALUE=19'b0000000_111000000001;
      15'b001_010011100101 : VALUE=19'b0000000_111000000000;
      15'b001_010011100110 : VALUE=19'b0000000_111000000000;
      15'b001_010011100111 : VALUE=19'b0000000_111000000000;
      15'b001_010011101000 : VALUE=19'b0000000_110111111111;
      15'b001_010011101001 : VALUE=19'b0000000_110111111111;
      15'b001_010011101010 : VALUE=19'b0000000_110111111111;
      15'b001_010011101011 : VALUE=19'b0000000_110111111110;
      15'b001_010011101100 : VALUE=19'b0000000_110111111110;
      15'b001_010011101101 : VALUE=19'b0000000_110111111110;
      15'b001_010011101110 : VALUE=19'b0000000_110111111101;
      15'b001_010011101111 : VALUE=19'b0000000_110111111101;
      15'b001_010011110000 : VALUE=19'b0000000_110111111101;
      15'b001_010011110001 : VALUE=19'b0000000_110111111100;
      15'b001_010011110010 : VALUE=19'b0000000_110111111100;
      15'b001_010011110011 : VALUE=19'b0000000_110111111100;
      15'b001_010011110100 : VALUE=19'b0000000_110111111011;
      15'b001_010011110101 : VALUE=19'b0000000_110111111011;
      15'b001_010011110110 : VALUE=19'b0000000_110111111011;
      15'b001_010011110111 : VALUE=19'b0000000_110111111010;
      15'b001_010011111000 : VALUE=19'b0000000_110111111010;
      15'b001_010011111001 : VALUE=19'b0000000_110111111010;
      15'b001_010011111010 : VALUE=19'b0000000_110111111001;
      15'b001_010011111011 : VALUE=19'b0000000_110111111001;
      15'b001_010011111100 : VALUE=19'b0000000_110111111001;
      15'b001_010011111101 : VALUE=19'b0000000_110111111000;
      15'b001_010011111110 : VALUE=19'b0000000_110111111000;
      15'b001_010011111111 : VALUE=19'b0000000_110111111000;
      15'b001_010100000000 : VALUE=19'b0000000_110111110111;
      15'b001_010100000001 : VALUE=19'b0000000_110111110111;
      15'b001_010100000010 : VALUE=19'b0000000_110111110111;
      15'b001_010100000011 : VALUE=19'b0000000_110111110110;
      15'b001_010100000100 : VALUE=19'b0000000_110111110110;
      15'b001_010100000101 : VALUE=19'b0000000_110111110110;
      15'b001_010100000110 : VALUE=19'b0000000_110111110101;
      15'b001_010100000111 : VALUE=19'b0000000_110111110101;
      15'b001_010100001000 : VALUE=19'b0000000_110111110101;
      15'b001_010100001001 : VALUE=19'b0000000_110111110100;
      15'b001_010100001010 : VALUE=19'b0000000_110111110100;
      15'b001_010100001011 : VALUE=19'b0000000_110111110100;
      15'b001_010100001100 : VALUE=19'b0000000_110111110011;
      15'b001_010100001101 : VALUE=19'b0000000_110111110011;
      15'b001_010100001110 : VALUE=19'b0000000_110111110011;
      15'b001_010100001111 : VALUE=19'b0000000_110111110010;
      15'b001_010100010000 : VALUE=19'b0000000_110111110010;
      15'b001_010100010001 : VALUE=19'b0000000_110111110010;
      15'b001_010100010010 : VALUE=19'b0000000_110111110001;
      15'b001_010100010011 : VALUE=19'b0000000_110111110001;
      15'b001_010100010100 : VALUE=19'b0000000_110111110001;
      15'b001_010100010101 : VALUE=19'b0000000_110111110000;
      15'b001_010100010110 : VALUE=19'b0000000_110111110000;
      15'b001_010100010111 : VALUE=19'b0000000_110111110000;
      15'b001_010100011000 : VALUE=19'b0000000_110111101111;
      15'b001_010100011001 : VALUE=19'b0000000_110111101111;
      15'b001_010100011010 : VALUE=19'b0000000_110111101111;
      15'b001_010100011011 : VALUE=19'b0000000_110111101110;
      15'b001_010100011100 : VALUE=19'b0000000_110111101110;
      15'b001_010100011101 : VALUE=19'b0000000_110111101110;
      15'b001_010100011110 : VALUE=19'b0000000_110111101101;
      15'b001_010100011111 : VALUE=19'b0000000_110111101101;
      15'b001_010100100000 : VALUE=19'b0000000_110111101101;
      15'b001_010100100001 : VALUE=19'b0000000_110111101100;
      15'b001_010100100010 : VALUE=19'b0000000_110111101100;
      15'b001_010100100011 : VALUE=19'b0000000_110111101100;
      15'b001_010100100100 : VALUE=19'b0000000_110111101011;
      15'b001_010100100101 : VALUE=19'b0000000_110111101011;
      15'b001_010100100110 : VALUE=19'b0000000_110111101011;
      15'b001_010100100111 : VALUE=19'b0000000_110111101010;
      15'b001_010100101000 : VALUE=19'b0000000_110111101010;
      15'b001_010100101001 : VALUE=19'b0000000_110111101010;
      15'b001_010100101010 : VALUE=19'b0000000_110111101001;
      15'b001_010100101011 : VALUE=19'b0000000_110111101001;
      15'b001_010100101100 : VALUE=19'b0000000_110111101001;
      15'b001_010100101101 : VALUE=19'b0000000_110111101000;
      15'b001_010100101110 : VALUE=19'b0000000_110111101000;
      15'b001_010100101111 : VALUE=19'b0000000_110111101000;
      15'b001_010100110000 : VALUE=19'b0000000_110111100111;
      15'b001_010100110001 : VALUE=19'b0000000_110111100111;
      15'b001_010100110010 : VALUE=19'b0000000_110111100111;
      15'b001_010100110011 : VALUE=19'b0000000_110111100110;
      15'b001_010100110100 : VALUE=19'b0000000_110111100110;
      15'b001_010100110101 : VALUE=19'b0000000_110111100110;
      15'b001_010100110110 : VALUE=19'b0000000_110111100101;
      15'b001_010100110111 : VALUE=19'b0000000_110111100101;
      15'b001_010100111000 : VALUE=19'b0000000_110111100101;
      15'b001_010100111001 : VALUE=19'b0000000_110111100100;
      15'b001_010100111010 : VALUE=19'b0000000_110111100100;
      15'b001_010100111011 : VALUE=19'b0000000_110111100100;
      15'b001_010100111100 : VALUE=19'b0000000_110111100011;
      15'b001_010100111101 : VALUE=19'b0000000_110111100011;
      15'b001_010100111110 : VALUE=19'b0000000_110111100011;
      15'b001_010100111111 : VALUE=19'b0000000_110111100011;
      15'b001_010101000000 : VALUE=19'b0000000_110111100010;
      15'b001_010101000001 : VALUE=19'b0000000_110111100010;
      15'b001_010101000010 : VALUE=19'b0000000_110111100010;
      15'b001_010101000011 : VALUE=19'b0000000_110111100001;
      15'b001_010101000100 : VALUE=19'b0000000_110111100001;
      15'b001_010101000101 : VALUE=19'b0000000_110111100001;
      15'b001_010101000110 : VALUE=19'b0000000_110111100000;
      15'b001_010101000111 : VALUE=19'b0000000_110111100000;
      15'b001_010101001000 : VALUE=19'b0000000_110111100000;
      15'b001_010101001001 : VALUE=19'b0000000_110111011111;
      15'b001_010101001010 : VALUE=19'b0000000_110111011111;
      15'b001_010101001011 : VALUE=19'b0000000_110111011111;
      15'b001_010101001100 : VALUE=19'b0000000_110111011110;
      15'b001_010101001101 : VALUE=19'b0000000_110111011110;
      15'b001_010101001110 : VALUE=19'b0000000_110111011110;
      15'b001_010101001111 : VALUE=19'b0000000_110111011101;
      15'b001_010101010000 : VALUE=19'b0000000_110111011101;
      15'b001_010101010001 : VALUE=19'b0000000_110111011101;
      15'b001_010101010010 : VALUE=19'b0000000_110111011100;
      15'b001_010101010011 : VALUE=19'b0000000_110111011100;
      15'b001_010101010100 : VALUE=19'b0000000_110111011100;
      15'b001_010101010101 : VALUE=19'b0000000_110111011011;
      15'b001_010101010110 : VALUE=19'b0000000_110111011011;
      15'b001_010101010111 : VALUE=19'b0000000_110111011011;
      15'b001_010101011000 : VALUE=19'b0000000_110111011010;
      15'b001_010101011001 : VALUE=19'b0000000_110111011010;
      15'b001_010101011010 : VALUE=19'b0000000_110111011010;
      15'b001_010101011011 : VALUE=19'b0000000_110111011001;
      15'b001_010101011100 : VALUE=19'b0000000_110111011001;
      15'b001_010101011101 : VALUE=19'b0000000_110111011001;
      15'b001_010101011110 : VALUE=19'b0000000_110111011000;
      15'b001_010101011111 : VALUE=19'b0000000_110111011000;
      15'b001_010101100000 : VALUE=19'b0000000_110111011000;
      15'b001_010101100001 : VALUE=19'b0000000_110111010111;
      15'b001_010101100010 : VALUE=19'b0000000_110111010111;
      15'b001_010101100011 : VALUE=19'b0000000_110111010111;
      15'b001_010101100100 : VALUE=19'b0000000_110111010110;
      15'b001_010101100101 : VALUE=19'b0000000_110111010110;
      15'b001_010101100110 : VALUE=19'b0000000_110111010110;
      15'b001_010101100111 : VALUE=19'b0000000_110111010110;
      15'b001_010101101000 : VALUE=19'b0000000_110111010101;
      15'b001_010101101001 : VALUE=19'b0000000_110111010101;
      15'b001_010101101010 : VALUE=19'b0000000_110111010101;
      15'b001_010101101011 : VALUE=19'b0000000_110111010100;
      15'b001_010101101100 : VALUE=19'b0000000_110111010100;
      15'b001_010101101101 : VALUE=19'b0000000_110111010100;
      15'b001_010101101110 : VALUE=19'b0000000_110111010011;
      15'b001_010101101111 : VALUE=19'b0000000_110111010011;
      15'b001_010101110000 : VALUE=19'b0000000_110111010011;
      15'b001_010101110001 : VALUE=19'b0000000_110111010010;
      15'b001_010101110010 : VALUE=19'b0000000_110111010010;
      15'b001_010101110011 : VALUE=19'b0000000_110111010010;
      15'b001_010101110100 : VALUE=19'b0000000_110111010001;
      15'b001_010101110101 : VALUE=19'b0000000_110111010001;
      15'b001_010101110110 : VALUE=19'b0000000_110111010001;
      15'b001_010101110111 : VALUE=19'b0000000_110111010000;
      15'b001_010101111000 : VALUE=19'b0000000_110111010000;
      15'b001_010101111001 : VALUE=19'b0000000_110111010000;
      15'b001_010101111010 : VALUE=19'b0000000_110111001111;
      15'b001_010101111011 : VALUE=19'b0000000_110111001111;
      15'b001_010101111100 : VALUE=19'b0000000_110111001111;
      15'b001_010101111101 : VALUE=19'b0000000_110111001110;
      15'b001_010101111110 : VALUE=19'b0000000_110111001110;
      15'b001_010101111111 : VALUE=19'b0000000_110111001110;
      15'b001_010110000000 : VALUE=19'b0000000_110111001101;
      15'b001_010110000001 : VALUE=19'b0000000_110111001101;
      15'b001_010110000010 : VALUE=19'b0000000_110111001101;
      15'b001_010110000011 : VALUE=19'b0000000_110111001101;
      15'b001_010110000100 : VALUE=19'b0000000_110111001100;
      15'b001_010110000101 : VALUE=19'b0000000_110111001100;
      15'b001_010110000110 : VALUE=19'b0000000_110111001100;
      15'b001_010110000111 : VALUE=19'b0000000_110111001011;
      15'b001_010110001000 : VALUE=19'b0000000_110111001011;
      15'b001_010110001001 : VALUE=19'b0000000_110111001011;
      15'b001_010110001010 : VALUE=19'b0000000_110111001010;
      15'b001_010110001011 : VALUE=19'b0000000_110111001010;
      15'b001_010110001100 : VALUE=19'b0000000_110111001010;
      15'b001_010110001101 : VALUE=19'b0000000_110111001001;
      15'b001_010110001110 : VALUE=19'b0000000_110111001001;
      15'b001_010110001111 : VALUE=19'b0000000_110111001001;
      15'b001_010110010000 : VALUE=19'b0000000_110111001000;
      15'b001_010110010001 : VALUE=19'b0000000_110111001000;
      15'b001_010110010010 : VALUE=19'b0000000_110111001000;
      15'b001_010110010011 : VALUE=19'b0000000_110111000111;
      15'b001_010110010100 : VALUE=19'b0000000_110111000111;
      15'b001_010110010101 : VALUE=19'b0000000_110111000111;
      15'b001_010110010110 : VALUE=19'b0000000_110111000110;
      15'b001_010110010111 : VALUE=19'b0000000_110111000110;
      15'b001_010110011000 : VALUE=19'b0000000_110111000110;
      15'b001_010110011001 : VALUE=19'b0000000_110111000101;
      15'b001_010110011010 : VALUE=19'b0000000_110111000101;
      15'b001_010110011011 : VALUE=19'b0000000_110111000101;
      15'b001_010110011100 : VALUE=19'b0000000_110111000101;
      15'b001_010110011101 : VALUE=19'b0000000_110111000100;
      15'b001_010110011110 : VALUE=19'b0000000_110111000100;
      15'b001_010110011111 : VALUE=19'b0000000_110111000100;
      15'b001_010110100000 : VALUE=19'b0000000_110111000011;
      15'b001_010110100001 : VALUE=19'b0000000_110111000011;
      15'b001_010110100010 : VALUE=19'b0000000_110111000011;
      15'b001_010110100011 : VALUE=19'b0000000_110111000010;
      15'b001_010110100100 : VALUE=19'b0000000_110111000010;
      15'b001_010110100101 : VALUE=19'b0000000_110111000010;
      15'b001_010110100110 : VALUE=19'b0000000_110111000001;
      15'b001_010110100111 : VALUE=19'b0000000_110111000001;
      15'b001_010110101000 : VALUE=19'b0000000_110111000001;
      15'b001_010110101001 : VALUE=19'b0000000_110111000000;
      15'b001_010110101010 : VALUE=19'b0000000_110111000000;
      15'b001_010110101011 : VALUE=19'b0000000_110111000000;
      15'b001_010110101100 : VALUE=19'b0000000_110110111111;
      15'b001_010110101101 : VALUE=19'b0000000_110110111111;
      15'b001_010110101110 : VALUE=19'b0000000_110110111111;
      15'b001_010110101111 : VALUE=19'b0000000_110110111110;
      15'b001_010110110000 : VALUE=19'b0000000_110110111110;
      15'b001_010110110001 : VALUE=19'b0000000_110110111110;
      15'b001_010110110010 : VALUE=19'b0000000_110110111110;
      15'b001_010110110011 : VALUE=19'b0000000_110110111101;
      15'b001_010110110100 : VALUE=19'b0000000_110110111101;
      15'b001_010110110101 : VALUE=19'b0000000_110110111101;
      15'b001_010110110110 : VALUE=19'b0000000_110110111100;
      15'b001_010110110111 : VALUE=19'b0000000_110110111100;
      15'b001_010110111000 : VALUE=19'b0000000_110110111100;
      15'b001_010110111001 : VALUE=19'b0000000_110110111011;
      15'b001_010110111010 : VALUE=19'b0000000_110110111011;
      15'b001_010110111011 : VALUE=19'b0000000_110110111011;
      15'b001_010110111100 : VALUE=19'b0000000_110110111010;
      15'b001_010110111101 : VALUE=19'b0000000_110110111010;
      15'b001_010110111110 : VALUE=19'b0000000_110110111010;
      15'b001_010110111111 : VALUE=19'b0000000_110110111001;
      15'b001_010111000000 : VALUE=19'b0000000_110110111001;
      15'b001_010111000001 : VALUE=19'b0000000_110110111001;
      15'b001_010111000010 : VALUE=19'b0000000_110110111000;
      15'b001_010111000011 : VALUE=19'b0000000_110110111000;
      15'b001_010111000100 : VALUE=19'b0000000_110110111000;
      15'b001_010111000101 : VALUE=19'b0000000_110110111000;
      15'b001_010111000110 : VALUE=19'b0000000_110110110111;
      15'b001_010111000111 : VALUE=19'b0000000_110110110111;
      15'b001_010111001000 : VALUE=19'b0000000_110110110111;
      15'b001_010111001001 : VALUE=19'b0000000_110110110110;
      15'b001_010111001010 : VALUE=19'b0000000_110110110110;
      15'b001_010111001011 : VALUE=19'b0000000_110110110110;
      15'b001_010111001100 : VALUE=19'b0000000_110110110101;
      15'b001_010111001101 : VALUE=19'b0000000_110110110101;
      15'b001_010111001110 : VALUE=19'b0000000_110110110101;
      15'b001_010111001111 : VALUE=19'b0000000_110110110100;
      15'b001_010111010000 : VALUE=19'b0000000_110110110100;
      15'b001_010111010001 : VALUE=19'b0000000_110110110100;
      15'b001_010111010010 : VALUE=19'b0000000_110110110011;
      15'b001_010111010011 : VALUE=19'b0000000_110110110011;
      15'b001_010111010100 : VALUE=19'b0000000_110110110011;
      15'b001_010111010101 : VALUE=19'b0000000_110110110010;
      15'b001_010111010110 : VALUE=19'b0000000_110110110010;
      15'b001_010111010111 : VALUE=19'b0000000_110110110010;
      15'b001_010111011000 : VALUE=19'b0000000_110110110010;
      15'b001_010111011001 : VALUE=19'b0000000_110110110001;
      15'b001_010111011010 : VALUE=19'b0000000_110110110001;
      15'b001_010111011011 : VALUE=19'b0000000_110110110001;
      15'b001_010111011100 : VALUE=19'b0000000_110110110000;
      15'b001_010111011101 : VALUE=19'b0000000_110110110000;
      15'b001_010111011110 : VALUE=19'b0000000_110110110000;
      15'b001_010111011111 : VALUE=19'b0000000_110110101111;
      15'b001_010111100000 : VALUE=19'b0000000_110110101111;
      15'b001_010111100001 : VALUE=19'b0000000_110110101111;
      15'b001_010111100010 : VALUE=19'b0000000_110110101110;
      15'b001_010111100011 : VALUE=19'b0000000_110110101110;
      15'b001_010111100100 : VALUE=19'b0000000_110110101110;
      15'b001_010111100101 : VALUE=19'b0000000_110110101101;
      15'b001_010111100110 : VALUE=19'b0000000_110110101101;
      15'b001_010111100111 : VALUE=19'b0000000_110110101101;
      15'b001_010111101000 : VALUE=19'b0000000_110110101101;
      15'b001_010111101001 : VALUE=19'b0000000_110110101100;
      15'b001_010111101010 : VALUE=19'b0000000_110110101100;
      15'b001_010111101011 : VALUE=19'b0000000_110110101100;
      15'b001_010111101100 : VALUE=19'b0000000_110110101011;
      15'b001_010111101101 : VALUE=19'b0000000_110110101011;
      15'b001_010111101110 : VALUE=19'b0000000_110110101011;
      15'b001_010111101111 : VALUE=19'b0000000_110110101010;
      15'b001_010111110000 : VALUE=19'b0000000_110110101010;
      15'b001_010111110001 : VALUE=19'b0000000_110110101010;
      15'b001_010111110010 : VALUE=19'b0000000_110110101001;
      15'b001_010111110011 : VALUE=19'b0000000_110110101001;
      15'b001_010111110100 : VALUE=19'b0000000_110110101001;
      15'b001_010111110101 : VALUE=19'b0000000_110110101000;
      15'b001_010111110110 : VALUE=19'b0000000_110110101000;
      15'b001_010111110111 : VALUE=19'b0000000_110110101000;
      15'b001_010111111000 : VALUE=19'b0000000_110110101000;
      15'b001_010111111001 : VALUE=19'b0000000_110110100111;
      15'b001_010111111010 : VALUE=19'b0000000_110110100111;
      15'b001_010111111011 : VALUE=19'b0000000_110110100111;
      15'b001_010111111100 : VALUE=19'b0000000_110110100110;
      15'b001_010111111101 : VALUE=19'b0000000_110110100110;
      15'b001_010111111110 : VALUE=19'b0000000_110110100110;
      15'b001_010111111111 : VALUE=19'b0000000_110110100101;
      15'b001_011000000000 : VALUE=19'b0000000_110110100101;
      15'b001_011000000001 : VALUE=19'b0000000_110110100101;
      15'b001_011000000010 : VALUE=19'b0000000_110110100100;
      15'b001_011000000011 : VALUE=19'b0000000_110110100100;
      15'b001_011000000100 : VALUE=19'b0000000_110110100100;
      15'b001_011000000101 : VALUE=19'b0000000_110110100100;
      15'b001_011000000110 : VALUE=19'b0000000_110110100011;
      15'b001_011000000111 : VALUE=19'b0000000_110110100011;
      15'b001_011000001000 : VALUE=19'b0000000_110110100011;
      15'b001_011000001001 : VALUE=19'b0000000_110110100010;
      15'b001_011000001010 : VALUE=19'b0000000_110110100010;
      15'b001_011000001011 : VALUE=19'b0000000_110110100010;
      15'b001_011000001100 : VALUE=19'b0000000_110110100001;
      15'b001_011000001101 : VALUE=19'b0000000_110110100001;
      15'b001_011000001110 : VALUE=19'b0000000_110110100001;
      15'b001_011000001111 : VALUE=19'b0000000_110110100000;
      15'b001_011000010000 : VALUE=19'b0000000_110110100000;
      15'b001_011000010001 : VALUE=19'b0000000_110110100000;
      15'b001_011000010010 : VALUE=19'b0000000_110110100000;
      15'b001_011000010011 : VALUE=19'b0000000_110110011111;
      15'b001_011000010100 : VALUE=19'b0000000_110110011111;
      15'b001_011000010101 : VALUE=19'b0000000_110110011111;
      15'b001_011000010110 : VALUE=19'b0000000_110110011110;
      15'b001_011000010111 : VALUE=19'b0000000_110110011110;
      15'b001_011000011000 : VALUE=19'b0000000_110110011110;
      15'b001_011000011001 : VALUE=19'b0000000_110110011101;
      15'b001_011000011010 : VALUE=19'b0000000_110110011101;
      15'b001_011000011011 : VALUE=19'b0000000_110110011101;
      15'b001_011000011100 : VALUE=19'b0000000_110110011100;
      15'b001_011000011101 : VALUE=19'b0000000_110110011100;
      15'b001_011000011110 : VALUE=19'b0000000_110110011100;
      15'b001_011000011111 : VALUE=19'b0000000_110110011100;
      15'b001_011000100000 : VALUE=19'b0000000_110110011011;
      15'b001_011000100001 : VALUE=19'b0000000_110110011011;
      15'b001_011000100010 : VALUE=19'b0000000_110110011011;
      15'b001_011000100011 : VALUE=19'b0000000_110110011010;
      15'b001_011000100100 : VALUE=19'b0000000_110110011010;
      15'b001_011000100101 : VALUE=19'b0000000_110110011010;
      15'b001_011000100110 : VALUE=19'b0000000_110110011001;
      15'b001_011000100111 : VALUE=19'b0000000_110110011001;
      15'b001_011000101000 : VALUE=19'b0000000_110110011001;
      15'b001_011000101001 : VALUE=19'b0000000_110110011000;
      15'b001_011000101010 : VALUE=19'b0000000_110110011000;
      15'b001_011000101011 : VALUE=19'b0000000_110110011000;
      15'b001_011000101100 : VALUE=19'b0000000_110110011000;
      15'b001_011000101101 : VALUE=19'b0000000_110110010111;
      15'b001_011000101110 : VALUE=19'b0000000_110110010111;
      15'b001_011000101111 : VALUE=19'b0000000_110110010111;
      15'b001_011000110000 : VALUE=19'b0000000_110110010110;
      15'b001_011000110001 : VALUE=19'b0000000_110110010110;
      15'b001_011000110010 : VALUE=19'b0000000_110110010110;
      15'b001_011000110011 : VALUE=19'b0000000_110110010101;
      15'b001_011000110100 : VALUE=19'b0000000_110110010101;
      15'b001_011000110101 : VALUE=19'b0000000_110110010101;
      15'b001_011000110110 : VALUE=19'b0000000_110110010100;
      15'b001_011000110111 : VALUE=19'b0000000_110110010100;
      15'b001_011000111000 : VALUE=19'b0000000_110110010100;
      15'b001_011000111001 : VALUE=19'b0000000_110110010100;
      15'b001_011000111010 : VALUE=19'b0000000_110110010011;
      15'b001_011000111011 : VALUE=19'b0000000_110110010011;
      15'b001_011000111100 : VALUE=19'b0000000_110110010011;
      15'b001_011000111101 : VALUE=19'b0000000_110110010010;
      15'b001_011000111110 : VALUE=19'b0000000_110110010010;
      15'b001_011000111111 : VALUE=19'b0000000_110110010010;
      15'b001_011001000000 : VALUE=19'b0000000_110110010001;
      15'b001_011001000001 : VALUE=19'b0000000_110110010001;
      15'b001_011001000010 : VALUE=19'b0000000_110110010001;
      15'b001_011001000011 : VALUE=19'b0000000_110110010000;
      15'b001_011001000100 : VALUE=19'b0000000_110110010000;
      15'b001_011001000101 : VALUE=19'b0000000_110110010000;
      15'b001_011001000110 : VALUE=19'b0000000_110110010000;
      15'b001_011001000111 : VALUE=19'b0000000_110110001111;
      15'b001_011001001000 : VALUE=19'b0000000_110110001111;
      15'b001_011001001001 : VALUE=19'b0000000_110110001111;
      15'b001_011001001010 : VALUE=19'b0000000_110110001110;
      15'b001_011001001011 : VALUE=19'b0000000_110110001110;
      15'b001_011001001100 : VALUE=19'b0000000_110110001110;
      15'b001_011001001101 : VALUE=19'b0000000_110110001101;
      15'b001_011001001110 : VALUE=19'b0000000_110110001101;
      15'b001_011001001111 : VALUE=19'b0000000_110110001101;
      15'b001_011001010000 : VALUE=19'b0000000_110110001101;
      15'b001_011001010001 : VALUE=19'b0000000_110110001100;
      15'b001_011001010010 : VALUE=19'b0000000_110110001100;
      15'b001_011001010011 : VALUE=19'b0000000_110110001100;
      15'b001_011001010100 : VALUE=19'b0000000_110110001011;
      15'b001_011001010101 : VALUE=19'b0000000_110110001011;
      15'b001_011001010110 : VALUE=19'b0000000_110110001011;
      15'b001_011001010111 : VALUE=19'b0000000_110110001010;
      15'b001_011001011000 : VALUE=19'b0000000_110110001010;
      15'b001_011001011001 : VALUE=19'b0000000_110110001010;
      15'b001_011001011010 : VALUE=19'b0000000_110110001010;
      15'b001_011001011011 : VALUE=19'b0000000_110110001001;
      15'b001_011001011100 : VALUE=19'b0000000_110110001001;
      15'b001_011001011101 : VALUE=19'b0000000_110110001001;
      15'b001_011001011110 : VALUE=19'b0000000_110110001000;
      15'b001_011001011111 : VALUE=19'b0000000_110110001000;
      15'b001_011001100000 : VALUE=19'b0000000_110110001000;
      15'b001_011001100001 : VALUE=19'b0000000_110110000111;
      15'b001_011001100010 : VALUE=19'b0000000_110110000111;
      15'b001_011001100011 : VALUE=19'b0000000_110110000111;
      15'b001_011001100100 : VALUE=19'b0000000_110110000110;
      15'b001_011001100101 : VALUE=19'b0000000_110110000110;
      15'b001_011001100110 : VALUE=19'b0000000_110110000110;
      15'b001_011001100111 : VALUE=19'b0000000_110110000110;
      15'b001_011001101000 : VALUE=19'b0000000_110110000101;
      15'b001_011001101001 : VALUE=19'b0000000_110110000101;
      15'b001_011001101010 : VALUE=19'b0000000_110110000101;
      15'b001_011001101011 : VALUE=19'b0000000_110110000100;
      15'b001_011001101100 : VALUE=19'b0000000_110110000100;
      15'b001_011001101101 : VALUE=19'b0000000_110110000100;
      15'b001_011001101110 : VALUE=19'b0000000_110110000011;
      15'b001_011001101111 : VALUE=19'b0000000_110110000011;
      15'b001_011001110000 : VALUE=19'b0000000_110110000011;
      15'b001_011001110001 : VALUE=19'b0000000_110110000011;
      15'b001_011001110010 : VALUE=19'b0000000_110110000010;
      15'b001_011001110011 : VALUE=19'b0000000_110110000010;
      15'b001_011001110100 : VALUE=19'b0000000_110110000010;
      15'b001_011001110101 : VALUE=19'b0000000_110110000001;
      15'b001_011001110110 : VALUE=19'b0000000_110110000001;
      15'b001_011001110111 : VALUE=19'b0000000_110110000001;
      15'b001_011001111000 : VALUE=19'b0000000_110110000000;
      15'b001_011001111001 : VALUE=19'b0000000_110110000000;
      15'b001_011001111010 : VALUE=19'b0000000_110110000000;
      15'b001_011001111011 : VALUE=19'b0000000_110110000000;
      15'b001_011001111100 : VALUE=19'b0000000_110101111111;
      15'b001_011001111101 : VALUE=19'b0000000_110101111111;
      15'b001_011001111110 : VALUE=19'b0000000_110101111111;
      15'b001_011001111111 : VALUE=19'b0000000_110101111110;
      15'b001_011010000000 : VALUE=19'b0000000_110101111110;
      15'b001_011010000001 : VALUE=19'b0000000_110101111110;
      15'b001_011010000010 : VALUE=19'b0000000_110101111101;
      15'b001_011010000011 : VALUE=19'b0000000_110101111101;
      15'b001_011010000100 : VALUE=19'b0000000_110101111101;
      15'b001_011010000101 : VALUE=19'b0000000_110101111101;
      15'b001_011010000110 : VALUE=19'b0000000_110101111100;
      15'b001_011010000111 : VALUE=19'b0000000_110101111100;
      15'b001_011010001000 : VALUE=19'b0000000_110101111100;
      15'b001_011010001001 : VALUE=19'b0000000_110101111011;
      15'b001_011010001010 : VALUE=19'b0000000_110101111011;
      15'b001_011010001011 : VALUE=19'b0000000_110101111011;
      15'b001_011010001100 : VALUE=19'b0000000_110101111010;
      15'b001_011010001101 : VALUE=19'b0000000_110101111010;
      15'b001_011010001110 : VALUE=19'b0000000_110101111010;
      15'b001_011010001111 : VALUE=19'b0000000_110101111010;
      15'b001_011010010000 : VALUE=19'b0000000_110101111001;
      15'b001_011010010001 : VALUE=19'b0000000_110101111001;
      15'b001_011010010010 : VALUE=19'b0000000_110101111001;
      15'b001_011010010011 : VALUE=19'b0000000_110101111000;
      15'b001_011010010100 : VALUE=19'b0000000_110101111000;
      15'b001_011010010101 : VALUE=19'b0000000_110101111000;
      15'b001_011010010110 : VALUE=19'b0000000_110101110111;
      15'b001_011010010111 : VALUE=19'b0000000_110101110111;
      15'b001_011010011000 : VALUE=19'b0000000_110101110111;
      15'b001_011010011001 : VALUE=19'b0000000_110101110111;
      15'b001_011010011010 : VALUE=19'b0000000_110101110110;
      15'b001_011010011011 : VALUE=19'b0000000_110101110110;
      15'b001_011010011100 : VALUE=19'b0000000_110101110110;
      15'b001_011010011101 : VALUE=19'b0000000_110101110101;
      15'b001_011010011110 : VALUE=19'b0000000_110101110101;
      15'b001_011010011111 : VALUE=19'b0000000_110101110101;
      15'b001_011010100000 : VALUE=19'b0000000_110101110100;
      15'b001_011010100001 : VALUE=19'b0000000_110101110100;
      15'b001_011010100010 : VALUE=19'b0000000_110101110100;
      15'b001_011010100011 : VALUE=19'b0000000_110101110100;
      15'b001_011010100100 : VALUE=19'b0000000_110101110011;
      15'b001_011010100101 : VALUE=19'b0000000_110101110011;
      15'b001_011010100110 : VALUE=19'b0000000_110101110011;
      15'b001_011010100111 : VALUE=19'b0000000_110101110010;
      15'b001_011010101000 : VALUE=19'b0000000_110101110010;
      15'b001_011010101001 : VALUE=19'b0000000_110101110010;
      15'b001_011010101010 : VALUE=19'b0000000_110101110010;
      15'b001_011010101011 : VALUE=19'b0000000_110101110001;
      15'b001_011010101100 : VALUE=19'b0000000_110101110001;
      15'b001_011010101101 : VALUE=19'b0000000_110101110001;
      15'b001_011010101110 : VALUE=19'b0000000_110101110000;
      15'b001_011010101111 : VALUE=19'b0000000_110101110000;
      15'b001_011010110000 : VALUE=19'b0000000_110101110000;
      15'b001_011010110001 : VALUE=19'b0000000_110101101111;
      15'b001_011010110010 : VALUE=19'b0000000_110101101111;
      15'b001_011010110011 : VALUE=19'b0000000_110101101111;
      15'b001_011010110100 : VALUE=19'b0000000_110101101111;
      15'b001_011010110101 : VALUE=19'b0000000_110101101110;
      15'b001_011010110110 : VALUE=19'b0000000_110101101110;
      15'b001_011010110111 : VALUE=19'b0000000_110101101110;
      15'b001_011010111000 : VALUE=19'b0000000_110101101101;
      15'b001_011010111001 : VALUE=19'b0000000_110101101101;
      15'b001_011010111010 : VALUE=19'b0000000_110101101101;
      15'b001_011010111011 : VALUE=19'b0000000_110101101100;
      15'b001_011010111100 : VALUE=19'b0000000_110101101100;
      15'b001_011010111101 : VALUE=19'b0000000_110101101100;
      15'b001_011010111110 : VALUE=19'b0000000_110101101100;
      15'b001_011010111111 : VALUE=19'b0000000_110101101011;
      15'b001_011011000000 : VALUE=19'b0000000_110101101011;
      15'b001_011011000001 : VALUE=19'b0000000_110101101011;
      15'b001_011011000010 : VALUE=19'b0000000_110101101010;
      15'b001_011011000011 : VALUE=19'b0000000_110101101010;
      15'b001_011011000100 : VALUE=19'b0000000_110101101010;
      15'b001_011011000101 : VALUE=19'b0000000_110101101010;
      15'b001_011011000110 : VALUE=19'b0000000_110101101001;
      15'b001_011011000111 : VALUE=19'b0000000_110101101001;
      15'b001_011011001000 : VALUE=19'b0000000_110101101001;
      15'b001_011011001001 : VALUE=19'b0000000_110101101000;
      15'b001_011011001010 : VALUE=19'b0000000_110101101000;
      15'b001_011011001011 : VALUE=19'b0000000_110101101000;
      15'b001_011011001100 : VALUE=19'b0000000_110101100111;
      15'b001_011011001101 : VALUE=19'b0000000_110101100111;
      15'b001_011011001110 : VALUE=19'b0000000_110101100111;
      15'b001_011011001111 : VALUE=19'b0000000_110101100111;
      15'b001_011011010000 : VALUE=19'b0000000_110101100110;
      15'b001_011011010001 : VALUE=19'b0000000_110101100110;
      15'b001_011011010010 : VALUE=19'b0000000_110101100110;
      15'b001_011011010011 : VALUE=19'b0000000_110101100101;
      15'b001_011011010100 : VALUE=19'b0000000_110101100101;
      15'b001_011011010101 : VALUE=19'b0000000_110101100101;
      15'b001_011011010110 : VALUE=19'b0000000_110101100101;
      15'b001_011011010111 : VALUE=19'b0000000_110101100100;
      15'b001_011011011000 : VALUE=19'b0000000_110101100100;
      15'b001_011011011001 : VALUE=19'b0000000_110101100100;
      15'b001_011011011010 : VALUE=19'b0000000_110101100011;
      15'b001_011011011011 : VALUE=19'b0000000_110101100011;
      15'b001_011011011100 : VALUE=19'b0000000_110101100011;
      15'b001_011011011101 : VALUE=19'b0000000_110101100010;
      15'b001_011011011110 : VALUE=19'b0000000_110101100010;
      15'b001_011011011111 : VALUE=19'b0000000_110101100010;
      15'b001_011011100000 : VALUE=19'b0000000_110101100010;
      15'b001_011011100001 : VALUE=19'b0000000_110101100001;
      15'b001_011011100010 : VALUE=19'b0000000_110101100001;
      15'b001_011011100011 : VALUE=19'b0000000_110101100001;
      15'b001_011011100100 : VALUE=19'b0000000_110101100000;
      15'b001_011011100101 : VALUE=19'b0000000_110101100000;
      15'b001_011011100110 : VALUE=19'b0000000_110101100000;
      15'b001_011011100111 : VALUE=19'b0000000_110101100000;
      15'b001_011011101000 : VALUE=19'b0000000_110101011111;
      15'b001_011011101001 : VALUE=19'b0000000_110101011111;
      15'b001_011011101010 : VALUE=19'b0000000_110101011111;
      15'b001_011011101011 : VALUE=19'b0000000_110101011110;
      15'b001_011011101100 : VALUE=19'b0000000_110101011110;
      15'b001_011011101101 : VALUE=19'b0000000_110101011110;
      15'b001_011011101110 : VALUE=19'b0000000_110101011110;
      15'b001_011011101111 : VALUE=19'b0000000_110101011101;
      15'b001_011011110000 : VALUE=19'b0000000_110101011101;
      15'b001_011011110001 : VALUE=19'b0000000_110101011101;
      15'b001_011011110010 : VALUE=19'b0000000_110101011100;
      15'b001_011011110011 : VALUE=19'b0000000_110101011100;
      15'b001_011011110100 : VALUE=19'b0000000_110101011100;
      15'b001_011011110101 : VALUE=19'b0000000_110101011011;
      15'b001_011011110110 : VALUE=19'b0000000_110101011011;
      15'b001_011011110111 : VALUE=19'b0000000_110101011011;
      15'b001_011011111000 : VALUE=19'b0000000_110101011011;
      15'b001_011011111001 : VALUE=19'b0000000_110101011010;
      15'b001_011011111010 : VALUE=19'b0000000_110101011010;
      15'b001_011011111011 : VALUE=19'b0000000_110101011010;
      15'b001_011011111100 : VALUE=19'b0000000_110101011001;
      15'b001_011011111101 : VALUE=19'b0000000_110101011001;
      15'b001_011011111110 : VALUE=19'b0000000_110101011001;
      15'b001_011011111111 : VALUE=19'b0000000_110101011001;
      15'b001_011100000000 : VALUE=19'b0000000_110101011000;
      15'b001_011100000001 : VALUE=19'b0000000_110101011000;
      15'b001_011100000010 : VALUE=19'b0000000_110101011000;
      15'b001_011100000011 : VALUE=19'b0000000_110101010111;
      15'b001_011100000100 : VALUE=19'b0000000_110101010111;
      15'b001_011100000101 : VALUE=19'b0000000_110101010111;
      15'b001_011100000110 : VALUE=19'b0000000_110101010111;
      15'b001_011100000111 : VALUE=19'b0000000_110101010110;
      15'b001_011100001000 : VALUE=19'b0000000_110101010110;
      15'b001_011100001001 : VALUE=19'b0000000_110101010110;
      15'b001_011100001010 : VALUE=19'b0000000_110101010101;
      15'b001_011100001011 : VALUE=19'b0000000_110101010101;
      15'b001_011100001100 : VALUE=19'b0000000_110101010101;
      15'b001_011100001101 : VALUE=19'b0000000_110101010101;
      15'b001_011100001110 : VALUE=19'b0000000_110101010100;
      15'b001_011100001111 : VALUE=19'b0000000_110101010100;
      15'b001_011100010000 : VALUE=19'b0000000_110101010100;
      15'b001_011100010001 : VALUE=19'b0000000_110101010011;
      15'b001_011100010010 : VALUE=19'b0000000_110101010011;
      15'b001_011100010011 : VALUE=19'b0000000_110101010011;
      15'b001_011100010100 : VALUE=19'b0000000_110101010011;
      15'b001_011100010101 : VALUE=19'b0000000_110101010010;
      15'b001_011100010110 : VALUE=19'b0000000_110101010010;
      15'b001_011100010111 : VALUE=19'b0000000_110101010010;
      15'b001_011100011000 : VALUE=19'b0000000_110101010001;
      15'b001_011100011001 : VALUE=19'b0000000_110101010001;
      15'b001_011100011010 : VALUE=19'b0000000_110101010001;
      15'b001_011100011011 : VALUE=19'b0000000_110101010000;
      15'b001_011100011100 : VALUE=19'b0000000_110101010000;
      15'b001_011100011101 : VALUE=19'b0000000_110101010000;
      15'b001_011100011110 : VALUE=19'b0000000_110101010000;
      15'b001_011100011111 : VALUE=19'b0000000_110101001111;
      15'b001_011100100000 : VALUE=19'b0000000_110101001111;
      15'b001_011100100001 : VALUE=19'b0000000_110101001111;
      15'b001_011100100010 : VALUE=19'b0000000_110101001110;
      15'b001_011100100011 : VALUE=19'b0000000_110101001110;
      15'b001_011100100100 : VALUE=19'b0000000_110101001110;
      15'b001_011100100101 : VALUE=19'b0000000_110101001110;
      15'b001_011100100110 : VALUE=19'b0000000_110101001101;
      15'b001_011100100111 : VALUE=19'b0000000_110101001101;
      15'b001_011100101000 : VALUE=19'b0000000_110101001101;
      15'b001_011100101001 : VALUE=19'b0000000_110101001100;
      15'b001_011100101010 : VALUE=19'b0000000_110101001100;
      15'b001_011100101011 : VALUE=19'b0000000_110101001100;
      15'b001_011100101100 : VALUE=19'b0000000_110101001100;
      15'b001_011100101101 : VALUE=19'b0000000_110101001011;
      15'b001_011100101110 : VALUE=19'b0000000_110101001011;
      15'b001_011100101111 : VALUE=19'b0000000_110101001011;
      15'b001_011100110000 : VALUE=19'b0000000_110101001010;
      15'b001_011100110001 : VALUE=19'b0000000_110101001010;
      15'b001_011100110010 : VALUE=19'b0000000_110101001010;
      15'b001_011100110011 : VALUE=19'b0000000_110101001010;
      15'b001_011100110100 : VALUE=19'b0000000_110101001001;
      15'b001_011100110101 : VALUE=19'b0000000_110101001001;
      15'b001_011100110110 : VALUE=19'b0000000_110101001001;
      15'b001_011100110111 : VALUE=19'b0000000_110101001000;
      15'b001_011100111000 : VALUE=19'b0000000_110101001000;
      15'b001_011100111001 : VALUE=19'b0000000_110101001000;
      15'b001_011100111010 : VALUE=19'b0000000_110101001000;
      15'b001_011100111011 : VALUE=19'b0000000_110101000111;
      15'b001_011100111100 : VALUE=19'b0000000_110101000111;
      15'b001_011100111101 : VALUE=19'b0000000_110101000111;
      15'b001_011100111110 : VALUE=19'b0000000_110101000110;
      15'b001_011100111111 : VALUE=19'b0000000_110101000110;
      15'b001_011101000000 : VALUE=19'b0000000_110101000110;
      15'b001_011101000001 : VALUE=19'b0000000_110101000110;
      15'b001_011101000010 : VALUE=19'b0000000_110101000101;
      15'b001_011101000011 : VALUE=19'b0000000_110101000101;
      15'b001_011101000100 : VALUE=19'b0000000_110101000101;
      15'b001_011101000101 : VALUE=19'b0000000_110101000100;
      15'b001_011101000110 : VALUE=19'b0000000_110101000100;
      15'b001_011101000111 : VALUE=19'b0000000_110101000100;
      15'b001_011101001000 : VALUE=19'b0000000_110101000100;
      15'b001_011101001001 : VALUE=19'b0000000_110101000011;
      15'b001_011101001010 : VALUE=19'b0000000_110101000011;
      15'b001_011101001011 : VALUE=19'b0000000_110101000011;
      15'b001_011101001100 : VALUE=19'b0000000_110101000010;
      15'b001_011101001101 : VALUE=19'b0000000_110101000010;
      15'b001_011101001110 : VALUE=19'b0000000_110101000010;
      15'b001_011101001111 : VALUE=19'b0000000_110101000010;
      15'b001_011101010000 : VALUE=19'b0000000_110101000001;
      15'b001_011101010001 : VALUE=19'b0000000_110101000001;
      15'b001_011101010010 : VALUE=19'b0000000_110101000001;
      15'b001_011101010011 : VALUE=19'b0000000_110101000000;
      15'b001_011101010100 : VALUE=19'b0000000_110101000000;
      15'b001_011101010101 : VALUE=19'b0000000_110101000000;
      15'b001_011101010110 : VALUE=19'b0000000_110101000000;
      15'b001_011101010111 : VALUE=19'b0000000_110100111111;
      15'b001_011101011000 : VALUE=19'b0000000_110100111111;
      15'b001_011101011001 : VALUE=19'b0000000_110100111111;
      15'b001_011101011010 : VALUE=19'b0000000_110100111110;
      15'b001_011101011011 : VALUE=19'b0000000_110100111110;
      15'b001_011101011100 : VALUE=19'b0000000_110100111110;
      15'b001_011101011101 : VALUE=19'b0000000_110100111110;
      15'b001_011101011110 : VALUE=19'b0000000_110100111101;
      15'b001_011101011111 : VALUE=19'b0000000_110100111101;
      15'b001_011101100000 : VALUE=19'b0000000_110100111101;
      15'b001_011101100001 : VALUE=19'b0000000_110100111101;
      15'b001_011101100010 : VALUE=19'b0000000_110100111100;
      15'b001_011101100011 : VALUE=19'b0000000_110100111100;
      15'b001_011101100100 : VALUE=19'b0000000_110100111100;
      15'b001_011101100101 : VALUE=19'b0000000_110100111011;
      15'b001_011101100110 : VALUE=19'b0000000_110100111011;
      15'b001_011101100111 : VALUE=19'b0000000_110100111011;
      15'b001_011101101000 : VALUE=19'b0000000_110100111011;
      15'b001_011101101001 : VALUE=19'b0000000_110100111010;
      15'b001_011101101010 : VALUE=19'b0000000_110100111010;
      15'b001_011101101011 : VALUE=19'b0000000_110100111010;
      15'b001_011101101100 : VALUE=19'b0000000_110100111001;
      15'b001_011101101101 : VALUE=19'b0000000_110100111001;
      15'b001_011101101110 : VALUE=19'b0000000_110100111001;
      15'b001_011101101111 : VALUE=19'b0000000_110100111001;
      15'b001_011101110000 : VALUE=19'b0000000_110100111000;
      15'b001_011101110001 : VALUE=19'b0000000_110100111000;
      15'b001_011101110010 : VALUE=19'b0000000_110100111000;
      15'b001_011101110011 : VALUE=19'b0000000_110100110111;
      15'b001_011101110100 : VALUE=19'b0000000_110100110111;
      15'b001_011101110101 : VALUE=19'b0000000_110100110111;
      15'b001_011101110110 : VALUE=19'b0000000_110100110111;
      15'b001_011101110111 : VALUE=19'b0000000_110100110110;
      15'b001_011101111000 : VALUE=19'b0000000_110100110110;
      15'b001_011101111001 : VALUE=19'b0000000_110100110110;
      15'b001_011101111010 : VALUE=19'b0000000_110100110101;
      15'b001_011101111011 : VALUE=19'b0000000_110100110101;
      15'b001_011101111100 : VALUE=19'b0000000_110100110101;
      15'b001_011101111101 : VALUE=19'b0000000_110100110101;
      15'b001_011101111110 : VALUE=19'b0000000_110100110100;
      15'b001_011101111111 : VALUE=19'b0000000_110100110100;
      15'b001_011110000000 : VALUE=19'b0000000_110100110100;
      15'b001_011110000001 : VALUE=19'b0000000_110100110011;
      15'b001_011110000010 : VALUE=19'b0000000_110100110011;
      15'b001_011110000011 : VALUE=19'b0000000_110100110011;
      15'b001_011110000100 : VALUE=19'b0000000_110100110011;
      15'b001_011110000101 : VALUE=19'b0000000_110100110010;
      15'b001_011110000110 : VALUE=19'b0000000_110100110010;
      15'b001_011110000111 : VALUE=19'b0000000_110100110010;
      15'b001_011110001000 : VALUE=19'b0000000_110100110010;
      15'b001_011110001001 : VALUE=19'b0000000_110100110001;
      15'b001_011110001010 : VALUE=19'b0000000_110100110001;
      15'b001_011110001011 : VALUE=19'b0000000_110100110001;
      15'b001_011110001100 : VALUE=19'b0000000_110100110000;
      15'b001_011110001101 : VALUE=19'b0000000_110100110000;
      15'b001_011110001110 : VALUE=19'b0000000_110100110000;
      15'b001_011110001111 : VALUE=19'b0000000_110100110000;
      15'b001_011110010000 : VALUE=19'b0000000_110100101111;
      15'b001_011110010001 : VALUE=19'b0000000_110100101111;
      15'b001_011110010010 : VALUE=19'b0000000_110100101111;
      15'b001_011110010011 : VALUE=19'b0000000_110100101110;
      15'b001_011110010100 : VALUE=19'b0000000_110100101110;
      15'b001_011110010101 : VALUE=19'b0000000_110100101110;
      15'b001_011110010110 : VALUE=19'b0000000_110100101110;
      15'b001_011110010111 : VALUE=19'b0000000_110100101101;
      15'b001_011110011000 : VALUE=19'b0000000_110100101101;
      15'b001_011110011001 : VALUE=19'b0000000_110100101101;
      15'b001_011110011010 : VALUE=19'b0000000_110100101100;
      15'b001_011110011011 : VALUE=19'b0000000_110100101100;
      15'b001_011110011100 : VALUE=19'b0000000_110100101100;
      15'b001_011110011101 : VALUE=19'b0000000_110100101100;
      15'b001_011110011110 : VALUE=19'b0000000_110100101011;
      15'b001_011110011111 : VALUE=19'b0000000_110100101011;
      15'b001_011110100000 : VALUE=19'b0000000_110100101011;
      15'b001_011110100001 : VALUE=19'b0000000_110100101011;
      15'b001_011110100010 : VALUE=19'b0000000_110100101010;
      15'b001_011110100011 : VALUE=19'b0000000_110100101010;
      15'b001_011110100100 : VALUE=19'b0000000_110100101010;
      15'b001_011110100101 : VALUE=19'b0000000_110100101001;
      15'b001_011110100110 : VALUE=19'b0000000_110100101001;
      15'b001_011110100111 : VALUE=19'b0000000_110100101001;
      15'b001_011110101000 : VALUE=19'b0000000_110100101001;
      15'b001_011110101001 : VALUE=19'b0000000_110100101000;
      15'b001_011110101010 : VALUE=19'b0000000_110100101000;
      15'b001_011110101011 : VALUE=19'b0000000_110100101000;
      15'b001_011110101100 : VALUE=19'b0000000_110100100111;
      15'b001_011110101101 : VALUE=19'b0000000_110100100111;
      15'b001_011110101110 : VALUE=19'b0000000_110100100111;
      15'b001_011110101111 : VALUE=19'b0000000_110100100111;
      15'b001_011110110000 : VALUE=19'b0000000_110100100110;
      15'b001_011110110001 : VALUE=19'b0000000_110100100110;
      15'b001_011110110010 : VALUE=19'b0000000_110100100110;
      15'b001_011110110011 : VALUE=19'b0000000_110100100110;
      15'b001_011110110100 : VALUE=19'b0000000_110100100101;
      15'b001_011110110101 : VALUE=19'b0000000_110100100101;
      15'b001_011110110110 : VALUE=19'b0000000_110100100101;
      15'b001_011110110111 : VALUE=19'b0000000_110100100100;
      15'b001_011110111000 : VALUE=19'b0000000_110100100100;
      15'b001_011110111001 : VALUE=19'b0000000_110100100100;
      15'b001_011110111010 : VALUE=19'b0000000_110100100100;
      15'b001_011110111011 : VALUE=19'b0000000_110100100011;
      15'b001_011110111100 : VALUE=19'b0000000_110100100011;
      15'b001_011110111101 : VALUE=19'b0000000_110100100011;
      15'b001_011110111110 : VALUE=19'b0000000_110100100010;
      15'b001_011110111111 : VALUE=19'b0000000_110100100010;
      15'b001_011111000000 : VALUE=19'b0000000_110100100010;
      15'b001_011111000001 : VALUE=19'b0000000_110100100010;
      15'b001_011111000010 : VALUE=19'b0000000_110100100001;
      15'b001_011111000011 : VALUE=19'b0000000_110100100001;
      15'b001_011111000100 : VALUE=19'b0000000_110100100001;
      15'b001_011111000101 : VALUE=19'b0000000_110100100001;
      15'b001_011111000110 : VALUE=19'b0000000_110100100000;
      15'b001_011111000111 : VALUE=19'b0000000_110100100000;
      15'b001_011111001000 : VALUE=19'b0000000_110100100000;
      15'b001_011111001001 : VALUE=19'b0000000_110100011111;
      15'b001_011111001010 : VALUE=19'b0000000_110100011111;
      15'b001_011111001011 : VALUE=19'b0000000_110100011111;
      15'b001_011111001100 : VALUE=19'b0000000_110100011111;
      15'b001_011111001101 : VALUE=19'b0000000_110100011110;
      15'b001_011111001110 : VALUE=19'b0000000_110100011110;
      15'b001_011111001111 : VALUE=19'b0000000_110100011110;
      15'b001_011111010000 : VALUE=19'b0000000_110100011110;
      15'b001_011111010001 : VALUE=19'b0000000_110100011101;
      15'b001_011111010010 : VALUE=19'b0000000_110100011101;
      15'b001_011111010011 : VALUE=19'b0000000_110100011101;
      15'b001_011111010100 : VALUE=19'b0000000_110100011100;
      15'b001_011111010101 : VALUE=19'b0000000_110100011100;
      15'b001_011111010110 : VALUE=19'b0000000_110100011100;
      15'b001_011111010111 : VALUE=19'b0000000_110100011100;
      15'b001_011111011000 : VALUE=19'b0000000_110100011011;
      15'b001_011111011001 : VALUE=19'b0000000_110100011011;
      15'b001_011111011010 : VALUE=19'b0000000_110100011011;
      15'b001_011111011011 : VALUE=19'b0000000_110100011010;
      15'b001_011111011100 : VALUE=19'b0000000_110100011010;
      15'b001_011111011101 : VALUE=19'b0000000_110100011010;
      15'b001_011111011110 : VALUE=19'b0000000_110100011010;
      15'b001_011111011111 : VALUE=19'b0000000_110100011001;
      15'b001_011111100000 : VALUE=19'b0000000_110100011001;
      15'b001_011111100001 : VALUE=19'b0000000_110100011001;
      15'b001_011111100010 : VALUE=19'b0000000_110100011001;
      15'b001_011111100011 : VALUE=19'b0000000_110100011000;
      15'b001_011111100100 : VALUE=19'b0000000_110100011000;
      15'b001_011111100101 : VALUE=19'b0000000_110100011000;
      15'b001_011111100110 : VALUE=19'b0000000_110100010111;
      15'b001_011111100111 : VALUE=19'b0000000_110100010111;
      15'b001_011111101000 : VALUE=19'b0000000_110100010111;
      15'b001_011111101001 : VALUE=19'b0000000_110100010111;
      15'b001_011111101010 : VALUE=19'b0000000_110100010110;
      15'b001_011111101011 : VALUE=19'b0000000_110100010110;
      15'b001_011111101100 : VALUE=19'b0000000_110100010110;
      15'b001_011111101101 : VALUE=19'b0000000_110100010110;
      15'b001_011111101110 : VALUE=19'b0000000_110100010101;
      15'b001_011111101111 : VALUE=19'b0000000_110100010101;
      15'b001_011111110000 : VALUE=19'b0000000_110100010101;
      15'b001_011111110001 : VALUE=19'b0000000_110100010100;
      15'b001_011111110010 : VALUE=19'b0000000_110100010100;
      15'b001_011111110011 : VALUE=19'b0000000_110100010100;
      15'b001_011111110100 : VALUE=19'b0000000_110100010100;
      15'b001_011111110101 : VALUE=19'b0000000_110100010011;
      15'b001_011111110110 : VALUE=19'b0000000_110100010011;
      15'b001_011111110111 : VALUE=19'b0000000_110100010011;
      15'b001_011111111000 : VALUE=19'b0000000_110100010011;
      15'b001_011111111001 : VALUE=19'b0000000_110100010010;
      15'b001_011111111010 : VALUE=19'b0000000_110100010010;
      15'b001_011111111011 : VALUE=19'b0000000_110100010010;
      15'b001_011111111100 : VALUE=19'b0000000_110100010001;
      15'b001_011111111101 : VALUE=19'b0000000_110100010001;
      15'b001_011111111110 : VALUE=19'b0000000_110100010001;
      15'b001_011111111111 : VALUE=19'b0000000_110100010001;
      15'b001_100000000000 : VALUE=19'b0000000_110100010000;
      15'b001_100000000001 : VALUE=19'b0000000_110100010000;
      15'b001_100000000010 : VALUE=19'b0000000_110100010000;
      15'b001_100000000011 : VALUE=19'b0000000_110100010000;
      15'b001_100000000100 : VALUE=19'b0000000_110100001111;
      15'b001_100000000101 : VALUE=19'b0000000_110100001111;
      15'b001_100000000110 : VALUE=19'b0000000_110100001111;
      15'b001_100000000111 : VALUE=19'b0000000_110100001110;
      15'b001_100000001000 : VALUE=19'b0000000_110100001110;
      15'b001_100000001001 : VALUE=19'b0000000_110100001110;
      15'b001_100000001010 : VALUE=19'b0000000_110100001110;
      15'b001_100000001011 : VALUE=19'b0000000_110100001101;
      15'b001_100000001100 : VALUE=19'b0000000_110100001101;
      15'b001_100000001101 : VALUE=19'b0000000_110100001101;
      15'b001_100000001110 : VALUE=19'b0000000_110100001101;
      15'b001_100000001111 : VALUE=19'b0000000_110100001100;
      15'b001_100000010000 : VALUE=19'b0000000_110100001100;
      15'b001_100000010001 : VALUE=19'b0000000_110100001100;
      15'b001_100000010010 : VALUE=19'b0000000_110100001011;
      15'b001_100000010011 : VALUE=19'b0000000_110100001011;
      15'b001_100000010100 : VALUE=19'b0000000_110100001011;
      15'b001_100000010101 : VALUE=19'b0000000_110100001011;
      15'b001_100000010110 : VALUE=19'b0000000_110100001010;
      15'b001_100000010111 : VALUE=19'b0000000_110100001010;
      15'b001_100000011000 : VALUE=19'b0000000_110100001010;
      15'b001_100000011001 : VALUE=19'b0000000_110100001010;
      15'b001_100000011010 : VALUE=19'b0000000_110100001001;
      15'b001_100000011011 : VALUE=19'b0000000_110100001001;
      15'b001_100000011100 : VALUE=19'b0000000_110100001001;
      15'b001_100000011101 : VALUE=19'b0000000_110100001001;
      15'b001_100000011110 : VALUE=19'b0000000_110100001000;
      15'b001_100000011111 : VALUE=19'b0000000_110100001000;
      15'b001_100000100000 : VALUE=19'b0000000_110100001000;
      15'b001_100000100001 : VALUE=19'b0000000_110100000111;
      15'b001_100000100010 : VALUE=19'b0000000_110100000111;
      15'b001_100000100011 : VALUE=19'b0000000_110100000111;
      15'b001_100000100100 : VALUE=19'b0000000_110100000111;
      15'b001_100000100101 : VALUE=19'b0000000_110100000110;
      15'b001_100000100110 : VALUE=19'b0000000_110100000110;
      15'b001_100000100111 : VALUE=19'b0000000_110100000110;
      15'b001_100000101000 : VALUE=19'b0000000_110100000110;
      15'b001_100000101001 : VALUE=19'b0000000_110100000101;
      15'b001_100000101010 : VALUE=19'b0000000_110100000101;
      15'b001_100000101011 : VALUE=19'b0000000_110100000101;
      15'b001_100000101100 : VALUE=19'b0000000_110100000100;
      15'b001_100000101101 : VALUE=19'b0000000_110100000100;
      15'b001_100000101110 : VALUE=19'b0000000_110100000100;
      15'b001_100000101111 : VALUE=19'b0000000_110100000100;
      15'b001_100000110000 : VALUE=19'b0000000_110100000011;
      15'b001_100000110001 : VALUE=19'b0000000_110100000011;
      15'b001_100000110010 : VALUE=19'b0000000_110100000011;
      15'b001_100000110011 : VALUE=19'b0000000_110100000011;
      15'b001_100000110100 : VALUE=19'b0000000_110100000010;
      15'b001_100000110101 : VALUE=19'b0000000_110100000010;
      15'b001_100000110110 : VALUE=19'b0000000_110100000010;
      15'b001_100000110111 : VALUE=19'b0000000_110100000010;
      15'b001_100000111000 : VALUE=19'b0000000_110100000001;
      15'b001_100000111001 : VALUE=19'b0000000_110100000001;
      15'b001_100000111010 : VALUE=19'b0000000_110100000001;
      15'b001_100000111011 : VALUE=19'b0000000_110100000000;
      15'b001_100000111100 : VALUE=19'b0000000_110100000000;
      15'b001_100000111101 : VALUE=19'b0000000_110100000000;
      15'b001_100000111110 : VALUE=19'b0000000_110100000000;
      15'b001_100000111111 : VALUE=19'b0000000_110011111111;
      15'b001_100001000000 : VALUE=19'b0000000_110011111111;
      15'b001_100001000001 : VALUE=19'b0000000_110011111111;
      15'b001_100001000010 : VALUE=19'b0000000_110011111111;
      15'b001_100001000011 : VALUE=19'b0000000_110011111110;
      15'b001_100001000100 : VALUE=19'b0000000_110011111110;
      15'b001_100001000101 : VALUE=19'b0000000_110011111110;
      15'b001_100001000110 : VALUE=19'b0000000_110011111101;
      15'b001_100001000111 : VALUE=19'b0000000_110011111101;
      15'b001_100001001000 : VALUE=19'b0000000_110011111101;
      15'b001_100001001001 : VALUE=19'b0000000_110011111101;
      15'b001_100001001010 : VALUE=19'b0000000_110011111100;
      15'b001_100001001011 : VALUE=19'b0000000_110011111100;
      15'b001_100001001100 : VALUE=19'b0000000_110011111100;
      15'b001_100001001101 : VALUE=19'b0000000_110011111100;
      15'b001_100001001110 : VALUE=19'b0000000_110011111011;
      15'b001_100001001111 : VALUE=19'b0000000_110011111011;
      15'b001_100001010000 : VALUE=19'b0000000_110011111011;
      15'b001_100001010001 : VALUE=19'b0000000_110011111011;
      15'b001_100001010010 : VALUE=19'b0000000_110011111010;
      15'b001_100001010011 : VALUE=19'b0000000_110011111010;
      15'b001_100001010100 : VALUE=19'b0000000_110011111010;
      15'b001_100001010101 : VALUE=19'b0000000_110011111001;
      15'b001_100001010110 : VALUE=19'b0000000_110011111001;
      15'b001_100001010111 : VALUE=19'b0000000_110011111001;
      15'b001_100001011000 : VALUE=19'b0000000_110011111001;
      15'b001_100001011001 : VALUE=19'b0000000_110011111000;
      15'b001_100001011010 : VALUE=19'b0000000_110011111000;
      15'b001_100001011011 : VALUE=19'b0000000_110011111000;
      15'b001_100001011100 : VALUE=19'b0000000_110011111000;
      15'b001_100001011101 : VALUE=19'b0000000_110011110111;
      15'b001_100001011110 : VALUE=19'b0000000_110011110111;
      15'b001_100001011111 : VALUE=19'b0000000_110011110111;
      15'b001_100001100000 : VALUE=19'b0000000_110011110111;
      15'b001_100001100001 : VALUE=19'b0000000_110011110110;
      15'b001_100001100010 : VALUE=19'b0000000_110011110110;
      15'b001_100001100011 : VALUE=19'b0000000_110011110110;
      15'b001_100001100100 : VALUE=19'b0000000_110011110101;
      15'b001_100001100101 : VALUE=19'b0000000_110011110101;
      15'b001_100001100110 : VALUE=19'b0000000_110011110101;
      15'b001_100001100111 : VALUE=19'b0000000_110011110101;
      15'b001_100001101000 : VALUE=19'b0000000_110011110100;
      15'b001_100001101001 : VALUE=19'b0000000_110011110100;
      15'b001_100001101010 : VALUE=19'b0000000_110011110100;
      15'b001_100001101011 : VALUE=19'b0000000_110011110100;
      15'b001_100001101100 : VALUE=19'b0000000_110011110011;
      15'b001_100001101101 : VALUE=19'b0000000_110011110011;
      15'b001_100001101110 : VALUE=19'b0000000_110011110011;
      15'b001_100001101111 : VALUE=19'b0000000_110011110011;
      15'b001_100001110000 : VALUE=19'b0000000_110011110010;
      15'b001_100001110001 : VALUE=19'b0000000_110011110010;
      15'b001_100001110010 : VALUE=19'b0000000_110011110010;
      15'b001_100001110011 : VALUE=19'b0000000_110011110010;
      15'b001_100001110100 : VALUE=19'b0000000_110011110001;
      15'b001_100001110101 : VALUE=19'b0000000_110011110001;
      15'b001_100001110110 : VALUE=19'b0000000_110011110001;
      15'b001_100001110111 : VALUE=19'b0000000_110011110000;
      15'b001_100001111000 : VALUE=19'b0000000_110011110000;
      15'b001_100001111001 : VALUE=19'b0000000_110011110000;
      15'b001_100001111010 : VALUE=19'b0000000_110011110000;
      15'b001_100001111011 : VALUE=19'b0000000_110011101111;
      15'b001_100001111100 : VALUE=19'b0000000_110011101111;
      15'b001_100001111101 : VALUE=19'b0000000_110011101111;
      15'b001_100001111110 : VALUE=19'b0000000_110011101111;
      15'b001_100001111111 : VALUE=19'b0000000_110011101110;
      15'b001_100010000000 : VALUE=19'b0000000_110011101110;
      15'b001_100010000001 : VALUE=19'b0000000_110011101110;
      15'b001_100010000010 : VALUE=19'b0000000_110011101110;
      15'b001_100010000011 : VALUE=19'b0000000_110011101101;
      15'b001_100010000100 : VALUE=19'b0000000_110011101101;
      15'b001_100010000101 : VALUE=19'b0000000_110011101101;
      15'b001_100010000110 : VALUE=19'b0000000_110011101100;
      15'b001_100010000111 : VALUE=19'b0000000_110011101100;
      15'b001_100010001000 : VALUE=19'b0000000_110011101100;
      15'b001_100010001001 : VALUE=19'b0000000_110011101100;
      15'b001_100010001010 : VALUE=19'b0000000_110011101011;
      15'b001_100010001011 : VALUE=19'b0000000_110011101011;
      15'b001_100010001100 : VALUE=19'b0000000_110011101011;
      15'b001_100010001101 : VALUE=19'b0000000_110011101011;
      15'b001_100010001110 : VALUE=19'b0000000_110011101010;
      15'b001_100010001111 : VALUE=19'b0000000_110011101010;
      15'b001_100010010000 : VALUE=19'b0000000_110011101010;
      15'b001_100010010001 : VALUE=19'b0000000_110011101010;
      15'b001_100010010010 : VALUE=19'b0000000_110011101001;
      15'b001_100010010011 : VALUE=19'b0000000_110011101001;
      15'b001_100010010100 : VALUE=19'b0000000_110011101001;
      15'b001_100010010101 : VALUE=19'b0000000_110011101001;
      15'b001_100010010110 : VALUE=19'b0000000_110011101000;
      15'b001_100010010111 : VALUE=19'b0000000_110011101000;
      15'b001_100010011000 : VALUE=19'b0000000_110011101000;
      15'b001_100010011001 : VALUE=19'b0000000_110011100111;
      15'b001_100010011010 : VALUE=19'b0000000_110011100111;
      15'b001_100010011011 : VALUE=19'b0000000_110011100111;
      15'b001_100010011100 : VALUE=19'b0000000_110011100111;
      15'b001_100010011101 : VALUE=19'b0000000_110011100110;
      15'b001_100010011110 : VALUE=19'b0000000_110011100110;
      15'b001_100010011111 : VALUE=19'b0000000_110011100110;
      15'b001_100010100000 : VALUE=19'b0000000_110011100110;
      15'b001_100010100001 : VALUE=19'b0000000_110011100101;
      15'b001_100010100010 : VALUE=19'b0000000_110011100101;
      15'b001_100010100011 : VALUE=19'b0000000_110011100101;
      15'b001_100010100100 : VALUE=19'b0000000_110011100101;
      15'b001_100010100101 : VALUE=19'b0000000_110011100100;
      15'b001_100010100110 : VALUE=19'b0000000_110011100100;
      15'b001_100010100111 : VALUE=19'b0000000_110011100100;
      15'b001_100010101000 : VALUE=19'b0000000_110011100100;
      15'b001_100010101001 : VALUE=19'b0000000_110011100011;
      15'b001_100010101010 : VALUE=19'b0000000_110011100011;
      15'b001_100010101011 : VALUE=19'b0000000_110011100011;
      15'b001_100010101100 : VALUE=19'b0000000_110011100011;
      15'b001_100010101101 : VALUE=19'b0000000_110011100010;
      15'b001_100010101110 : VALUE=19'b0000000_110011100010;
      15'b001_100010101111 : VALUE=19'b0000000_110011100010;
      15'b001_100010110000 : VALUE=19'b0000000_110011100001;
      15'b001_100010110001 : VALUE=19'b0000000_110011100001;
      15'b001_100010110010 : VALUE=19'b0000000_110011100001;
      15'b001_100010110011 : VALUE=19'b0000000_110011100001;
      15'b001_100010110100 : VALUE=19'b0000000_110011100000;
      15'b001_100010110101 : VALUE=19'b0000000_110011100000;
      15'b001_100010110110 : VALUE=19'b0000000_110011100000;
      15'b001_100010110111 : VALUE=19'b0000000_110011100000;
      15'b001_100010111000 : VALUE=19'b0000000_110011011111;
      15'b001_100010111001 : VALUE=19'b0000000_110011011111;
      15'b001_100010111010 : VALUE=19'b0000000_110011011111;
      15'b001_100010111011 : VALUE=19'b0000000_110011011111;
      15'b001_100010111100 : VALUE=19'b0000000_110011011110;
      15'b001_100010111101 : VALUE=19'b0000000_110011011110;
      15'b001_100010111110 : VALUE=19'b0000000_110011011110;
      15'b001_100010111111 : VALUE=19'b0000000_110011011110;
      15'b001_100011000000 : VALUE=19'b0000000_110011011101;
      15'b001_100011000001 : VALUE=19'b0000000_110011011101;
      15'b001_100011000010 : VALUE=19'b0000000_110011011101;
      15'b001_100011000011 : VALUE=19'b0000000_110011011101;
      15'b001_100011000100 : VALUE=19'b0000000_110011011100;
      15'b001_100011000101 : VALUE=19'b0000000_110011011100;
      15'b001_100011000110 : VALUE=19'b0000000_110011011100;
      15'b001_100011000111 : VALUE=19'b0000000_110011011011;
      15'b001_100011001000 : VALUE=19'b0000000_110011011011;
      15'b001_100011001001 : VALUE=19'b0000000_110011011011;
      15'b001_100011001010 : VALUE=19'b0000000_110011011011;
      15'b001_100011001011 : VALUE=19'b0000000_110011011010;
      15'b001_100011001100 : VALUE=19'b0000000_110011011010;
      15'b001_100011001101 : VALUE=19'b0000000_110011011010;
      15'b001_100011001110 : VALUE=19'b0000000_110011011010;
      15'b001_100011001111 : VALUE=19'b0000000_110011011001;
      15'b001_100011010000 : VALUE=19'b0000000_110011011001;
      15'b001_100011010001 : VALUE=19'b0000000_110011011001;
      15'b001_100011010010 : VALUE=19'b0000000_110011011001;
      15'b001_100011010011 : VALUE=19'b0000000_110011011000;
      15'b001_100011010100 : VALUE=19'b0000000_110011011000;
      15'b001_100011010101 : VALUE=19'b0000000_110011011000;
      15'b001_100011010110 : VALUE=19'b0000000_110011011000;
      15'b001_100011010111 : VALUE=19'b0000000_110011010111;
      15'b001_100011011000 : VALUE=19'b0000000_110011010111;
      15'b001_100011011001 : VALUE=19'b0000000_110011010111;
      15'b001_100011011010 : VALUE=19'b0000000_110011010111;
      15'b001_100011011011 : VALUE=19'b0000000_110011010110;
      15'b001_100011011100 : VALUE=19'b0000000_110011010110;
      15'b001_100011011101 : VALUE=19'b0000000_110011010110;
      15'b001_100011011110 : VALUE=19'b0000000_110011010110;
      15'b001_100011011111 : VALUE=19'b0000000_110011010101;
      15'b001_100011100000 : VALUE=19'b0000000_110011010101;
      15'b001_100011100001 : VALUE=19'b0000000_110011010101;
      15'b001_100011100010 : VALUE=19'b0000000_110011010101;
      15'b001_100011100011 : VALUE=19'b0000000_110011010100;
      15'b001_100011100100 : VALUE=19'b0000000_110011010100;
      15'b001_100011100101 : VALUE=19'b0000000_110011010100;
      15'b001_100011100110 : VALUE=19'b0000000_110011010011;
      15'b001_100011100111 : VALUE=19'b0000000_110011010011;
      15'b001_100011101000 : VALUE=19'b0000000_110011010011;
      15'b001_100011101001 : VALUE=19'b0000000_110011010011;
      15'b001_100011101010 : VALUE=19'b0000000_110011010010;
      15'b001_100011101011 : VALUE=19'b0000000_110011010010;
      15'b001_100011101100 : VALUE=19'b0000000_110011010010;
      15'b001_100011101101 : VALUE=19'b0000000_110011010010;
      15'b001_100011101110 : VALUE=19'b0000000_110011010001;
      15'b001_100011101111 : VALUE=19'b0000000_110011010001;
      15'b001_100011110000 : VALUE=19'b0000000_110011010001;
      15'b001_100011110001 : VALUE=19'b0000000_110011010001;
      15'b001_100011110010 : VALUE=19'b0000000_110011010000;
      15'b001_100011110011 : VALUE=19'b0000000_110011010000;
      15'b001_100011110100 : VALUE=19'b0000000_110011010000;
      15'b001_100011110101 : VALUE=19'b0000000_110011010000;
      15'b001_100011110110 : VALUE=19'b0000000_110011001111;
      15'b001_100011110111 : VALUE=19'b0000000_110011001111;
      15'b001_100011111000 : VALUE=19'b0000000_110011001111;
      15'b001_100011111001 : VALUE=19'b0000000_110011001111;
      15'b001_100011111010 : VALUE=19'b0000000_110011001110;
      15'b001_100011111011 : VALUE=19'b0000000_110011001110;
      15'b001_100011111100 : VALUE=19'b0000000_110011001110;
      15'b001_100011111101 : VALUE=19'b0000000_110011001110;
      15'b001_100011111110 : VALUE=19'b0000000_110011001101;
      15'b001_100011111111 : VALUE=19'b0000000_110011001101;
      15'b001_100100000000 : VALUE=19'b0000000_110011001101;
      15'b001_100100000001 : VALUE=19'b0000000_110011001101;
      15'b001_100100000010 : VALUE=19'b0000000_110011001100;
      15'b001_100100000011 : VALUE=19'b0000000_110011001100;
      15'b001_100100000100 : VALUE=19'b0000000_110011001100;
      15'b001_100100000101 : VALUE=19'b0000000_110011001100;
      15'b001_100100000110 : VALUE=19'b0000000_110011001011;
      15'b001_100100000111 : VALUE=19'b0000000_110011001011;
      15'b001_100100001000 : VALUE=19'b0000000_110011001011;
      15'b001_100100001001 : VALUE=19'b0000000_110011001010;
      15'b001_100100001010 : VALUE=19'b0000000_110011001010;
      15'b001_100100001011 : VALUE=19'b0000000_110011001010;
      15'b001_100100001100 : VALUE=19'b0000000_110011001010;
      15'b001_100100001101 : VALUE=19'b0000000_110011001001;
      15'b001_100100001110 : VALUE=19'b0000000_110011001001;
      15'b001_100100001111 : VALUE=19'b0000000_110011001001;
      15'b001_100100010000 : VALUE=19'b0000000_110011001001;
      15'b001_100100010001 : VALUE=19'b0000000_110011001000;
      15'b001_100100010010 : VALUE=19'b0000000_110011001000;
      15'b001_100100010011 : VALUE=19'b0000000_110011001000;
      15'b001_100100010100 : VALUE=19'b0000000_110011001000;
      15'b001_100100010101 : VALUE=19'b0000000_110011000111;
      15'b001_100100010110 : VALUE=19'b0000000_110011000111;
      15'b001_100100010111 : VALUE=19'b0000000_110011000111;
      15'b001_100100011000 : VALUE=19'b0000000_110011000111;
      15'b001_100100011001 : VALUE=19'b0000000_110011000110;
      15'b001_100100011010 : VALUE=19'b0000000_110011000110;
      15'b001_100100011011 : VALUE=19'b0000000_110011000110;
      15'b001_100100011100 : VALUE=19'b0000000_110011000110;
      15'b001_100100011101 : VALUE=19'b0000000_110011000101;
      15'b001_100100011110 : VALUE=19'b0000000_110011000101;
      15'b001_100100011111 : VALUE=19'b0000000_110011000101;
      15'b001_100100100000 : VALUE=19'b0000000_110011000101;
      15'b001_100100100001 : VALUE=19'b0000000_110011000100;
      15'b001_100100100010 : VALUE=19'b0000000_110011000100;
      15'b001_100100100011 : VALUE=19'b0000000_110011000100;
      15'b001_100100100100 : VALUE=19'b0000000_110011000100;
      15'b001_100100100101 : VALUE=19'b0000000_110011000011;
      15'b001_100100100110 : VALUE=19'b0000000_110011000011;
      15'b001_100100100111 : VALUE=19'b0000000_110011000011;
      15'b001_100100101000 : VALUE=19'b0000000_110011000011;
      15'b001_100100101001 : VALUE=19'b0000000_110011000010;
      15'b001_100100101010 : VALUE=19'b0000000_110011000010;
      15'b001_100100101011 : VALUE=19'b0000000_110011000010;
      15'b001_100100101100 : VALUE=19'b0000000_110011000010;
      15'b001_100100101101 : VALUE=19'b0000000_110011000001;
      15'b001_100100101110 : VALUE=19'b0000000_110011000001;
      15'b001_100100101111 : VALUE=19'b0000000_110011000001;
      15'b001_100100110000 : VALUE=19'b0000000_110011000001;
      15'b001_100100110001 : VALUE=19'b0000000_110011000000;
      15'b001_100100110010 : VALUE=19'b0000000_110011000000;
      15'b001_100100110011 : VALUE=19'b0000000_110011000000;
      15'b001_100100110100 : VALUE=19'b0000000_110011000000;
      15'b001_100100110101 : VALUE=19'b0000000_110010111111;
      15'b001_100100110110 : VALUE=19'b0000000_110010111111;
      15'b001_100100110111 : VALUE=19'b0000000_110010111111;
      15'b001_100100111000 : VALUE=19'b0000000_110010111111;
      15'b001_100100111001 : VALUE=19'b0000000_110010111110;
      15'b001_100100111010 : VALUE=19'b0000000_110010111110;
      15'b001_100100111011 : VALUE=19'b0000000_110010111110;
      15'b001_100100111100 : VALUE=19'b0000000_110010111110;
      15'b001_100100111101 : VALUE=19'b0000000_110010111101;
      15'b001_100100111110 : VALUE=19'b0000000_110010111101;
      15'b001_100100111111 : VALUE=19'b0000000_110010111101;
      15'b001_100101000000 : VALUE=19'b0000000_110010111101;
      15'b001_100101000001 : VALUE=19'b0000000_110010111100;
      15'b001_100101000010 : VALUE=19'b0000000_110010111100;
      15'b001_100101000011 : VALUE=19'b0000000_110010111100;
      15'b001_100101000100 : VALUE=19'b0000000_110010111100;
      15'b001_100101000101 : VALUE=19'b0000000_110010111011;
      15'b001_100101000110 : VALUE=19'b0000000_110010111011;
      15'b001_100101000111 : VALUE=19'b0000000_110010111011;
      15'b001_100101001000 : VALUE=19'b0000000_110010111011;
      15'b001_100101001001 : VALUE=19'b0000000_110010111010;
      15'b001_100101001010 : VALUE=19'b0000000_110010111010;
      15'b001_100101001011 : VALUE=19'b0000000_110010111010;
      15'b001_100101001100 : VALUE=19'b0000000_110010111010;
      15'b001_100101001101 : VALUE=19'b0000000_110010111001;
      15'b001_100101001110 : VALUE=19'b0000000_110010111001;
      15'b001_100101001111 : VALUE=19'b0000000_110010111001;
      15'b001_100101010000 : VALUE=19'b0000000_110010111001;
      15'b001_100101010001 : VALUE=19'b0000000_110010111000;
      15'b001_100101010010 : VALUE=19'b0000000_110010111000;
      15'b001_100101010011 : VALUE=19'b0000000_110010111000;
      15'b001_100101010100 : VALUE=19'b0000000_110010111000;
      15'b001_100101010101 : VALUE=19'b0000000_110010110111;
      15'b001_100101010110 : VALUE=19'b0000000_110010110111;
      15'b001_100101010111 : VALUE=19'b0000000_110010110111;
      15'b001_100101011000 : VALUE=19'b0000000_110010110111;
      15'b001_100101011001 : VALUE=19'b0000000_110010110110;
      15'b001_100101011010 : VALUE=19'b0000000_110010110110;
      15'b001_100101011011 : VALUE=19'b0000000_110010110110;
      15'b001_100101011100 : VALUE=19'b0000000_110010110101;
      15'b001_100101011101 : VALUE=19'b0000000_110010110101;
      15'b001_100101011110 : VALUE=19'b0000000_110010110101;
      15'b001_100101011111 : VALUE=19'b0000000_110010110101;
      15'b001_100101100000 : VALUE=19'b0000000_110010110100;
      15'b001_100101100001 : VALUE=19'b0000000_110010110100;
      15'b001_100101100010 : VALUE=19'b0000000_110010110100;
      15'b001_100101100011 : VALUE=19'b0000000_110010110100;
      15'b001_100101100100 : VALUE=19'b0000000_110010110011;
      15'b001_100101100101 : VALUE=19'b0000000_110010110011;
      15'b001_100101100110 : VALUE=19'b0000000_110010110011;
      15'b001_100101100111 : VALUE=19'b0000000_110010110011;
      15'b001_100101101000 : VALUE=19'b0000000_110010110010;
      15'b001_100101101001 : VALUE=19'b0000000_110010110010;
      15'b001_100101101010 : VALUE=19'b0000000_110010110010;
      15'b001_100101101011 : VALUE=19'b0000000_110010110010;
      15'b001_100101101100 : VALUE=19'b0000000_110010110001;
      15'b001_100101101101 : VALUE=19'b0000000_110010110001;
      15'b001_100101101110 : VALUE=19'b0000000_110010110001;
      15'b001_100101101111 : VALUE=19'b0000000_110010110001;
      15'b001_100101110000 : VALUE=19'b0000000_110010110000;
      15'b001_100101110001 : VALUE=19'b0000000_110010110000;
      15'b001_100101110010 : VALUE=19'b0000000_110010110000;
      15'b001_100101110011 : VALUE=19'b0000000_110010110000;
      15'b001_100101110100 : VALUE=19'b0000000_110010110000;
      15'b001_100101110101 : VALUE=19'b0000000_110010101111;
      15'b001_100101110110 : VALUE=19'b0000000_110010101111;
      15'b001_100101110111 : VALUE=19'b0000000_110010101111;
      15'b001_100101111000 : VALUE=19'b0000000_110010101111;
      15'b001_100101111001 : VALUE=19'b0000000_110010101110;
      15'b001_100101111010 : VALUE=19'b0000000_110010101110;
      15'b001_100101111011 : VALUE=19'b0000000_110010101110;
      15'b001_100101111100 : VALUE=19'b0000000_110010101110;
      15'b001_100101111101 : VALUE=19'b0000000_110010101101;
      15'b001_100101111110 : VALUE=19'b0000000_110010101101;
      15'b001_100101111111 : VALUE=19'b0000000_110010101101;
      15'b001_100110000000 : VALUE=19'b0000000_110010101101;
      15'b001_100110000001 : VALUE=19'b0000000_110010101100;
      15'b001_100110000010 : VALUE=19'b0000000_110010101100;
      15'b001_100110000011 : VALUE=19'b0000000_110010101100;
      15'b001_100110000100 : VALUE=19'b0000000_110010101100;
      15'b001_100110000101 : VALUE=19'b0000000_110010101011;
      15'b001_100110000110 : VALUE=19'b0000000_110010101011;
      15'b001_100110000111 : VALUE=19'b0000000_110010101011;
      15'b001_100110001000 : VALUE=19'b0000000_110010101011;
      15'b001_100110001001 : VALUE=19'b0000000_110010101010;
      15'b001_100110001010 : VALUE=19'b0000000_110010101010;
      15'b001_100110001011 : VALUE=19'b0000000_110010101010;
      15'b001_100110001100 : VALUE=19'b0000000_110010101010;
      15'b001_100110001101 : VALUE=19'b0000000_110010101001;
      15'b001_100110001110 : VALUE=19'b0000000_110010101001;
      15'b001_100110001111 : VALUE=19'b0000000_110010101001;
      15'b001_100110010000 : VALUE=19'b0000000_110010101001;
      15'b001_100110010001 : VALUE=19'b0000000_110010101000;
      15'b001_100110010010 : VALUE=19'b0000000_110010101000;
      15'b001_100110010011 : VALUE=19'b0000000_110010101000;
      15'b001_100110010100 : VALUE=19'b0000000_110010101000;
      15'b001_100110010101 : VALUE=19'b0000000_110010100111;
      15'b001_100110010110 : VALUE=19'b0000000_110010100111;
      15'b001_100110010111 : VALUE=19'b0000000_110010100111;
      15'b001_100110011000 : VALUE=19'b0000000_110010100111;
      15'b001_100110011001 : VALUE=19'b0000000_110010100110;
      15'b001_100110011010 : VALUE=19'b0000000_110010100110;
      15'b001_100110011011 : VALUE=19'b0000000_110010100110;
      15'b001_100110011100 : VALUE=19'b0000000_110010100110;
      15'b001_100110011101 : VALUE=19'b0000000_110010100101;
      15'b001_100110011110 : VALUE=19'b0000000_110010100101;
      15'b001_100110011111 : VALUE=19'b0000000_110010100101;
      15'b001_100110100000 : VALUE=19'b0000000_110010100101;
      15'b001_100110100001 : VALUE=19'b0000000_110010100100;
      15'b001_100110100010 : VALUE=19'b0000000_110010100100;
      15'b001_100110100011 : VALUE=19'b0000000_110010100100;
      15'b001_100110100100 : VALUE=19'b0000000_110010100100;
      15'b001_100110100101 : VALUE=19'b0000000_110010100011;
      15'b001_100110100110 : VALUE=19'b0000000_110010100011;
      15'b001_100110100111 : VALUE=19'b0000000_110010100011;
      15'b001_100110101000 : VALUE=19'b0000000_110010100011;
      15'b001_100110101001 : VALUE=19'b0000000_110010100010;
      15'b001_100110101010 : VALUE=19'b0000000_110010100010;
      15'b001_100110101011 : VALUE=19'b0000000_110010100010;
      15'b001_100110101100 : VALUE=19'b0000000_110010100010;
      15'b001_100110101101 : VALUE=19'b0000000_110010100001;
      15'b001_100110101110 : VALUE=19'b0000000_110010100001;
      15'b001_100110101111 : VALUE=19'b0000000_110010100001;
      15'b001_100110110000 : VALUE=19'b0000000_110010100001;
      15'b001_100110110001 : VALUE=19'b0000000_110010100000;
      15'b001_100110110010 : VALUE=19'b0000000_110010100000;
      15'b001_100110110011 : VALUE=19'b0000000_110010100000;
      15'b001_100110110100 : VALUE=19'b0000000_110010100000;
      15'b001_100110110101 : VALUE=19'b0000000_110010011111;
      15'b001_100110110110 : VALUE=19'b0000000_110010011111;
      15'b001_100110110111 : VALUE=19'b0000000_110010011111;
      15'b001_100110111000 : VALUE=19'b0000000_110010011111;
      15'b001_100110111001 : VALUE=19'b0000000_110010011110;
      15'b001_100110111010 : VALUE=19'b0000000_110010011110;
      15'b001_100110111011 : VALUE=19'b0000000_110010011110;
      15'b001_100110111100 : VALUE=19'b0000000_110010011110;
      15'b001_100110111101 : VALUE=19'b0000000_110010011101;
      15'b001_100110111110 : VALUE=19'b0000000_110010011101;
      15'b001_100110111111 : VALUE=19'b0000000_110010011101;
      15'b001_100111000000 : VALUE=19'b0000000_110010011101;
      15'b001_100111000001 : VALUE=19'b0000000_110010011100;
      15'b001_100111000010 : VALUE=19'b0000000_110010011100;
      15'b001_100111000011 : VALUE=19'b0000000_110010011100;
      15'b001_100111000100 : VALUE=19'b0000000_110010011100;
      15'b001_100111000101 : VALUE=19'b0000000_110010011100;
      15'b001_100111000110 : VALUE=19'b0000000_110010011011;
      15'b001_100111000111 : VALUE=19'b0000000_110010011011;
      15'b001_100111001000 : VALUE=19'b0000000_110010011011;
      15'b001_100111001001 : VALUE=19'b0000000_110010011011;
      15'b001_100111001010 : VALUE=19'b0000000_110010011010;
      15'b001_100111001011 : VALUE=19'b0000000_110010011010;
      15'b001_100111001100 : VALUE=19'b0000000_110010011010;
      15'b001_100111001101 : VALUE=19'b0000000_110010011010;
      15'b001_100111001110 : VALUE=19'b0000000_110010011001;
      15'b001_100111001111 : VALUE=19'b0000000_110010011001;
      15'b001_100111010000 : VALUE=19'b0000000_110010011001;
      15'b001_100111010001 : VALUE=19'b0000000_110010011001;
      15'b001_100111010010 : VALUE=19'b0000000_110010011000;
      15'b001_100111010011 : VALUE=19'b0000000_110010011000;
      15'b001_100111010100 : VALUE=19'b0000000_110010011000;
      15'b001_100111010101 : VALUE=19'b0000000_110010011000;
      15'b001_100111010110 : VALUE=19'b0000000_110010010111;
      15'b001_100111010111 : VALUE=19'b0000000_110010010111;
      15'b001_100111011000 : VALUE=19'b0000000_110010010111;
      15'b001_100111011001 : VALUE=19'b0000000_110010010111;
      15'b001_100111011010 : VALUE=19'b0000000_110010010110;
      15'b001_100111011011 : VALUE=19'b0000000_110010010110;
      15'b001_100111011100 : VALUE=19'b0000000_110010010110;
      15'b001_100111011101 : VALUE=19'b0000000_110010010110;
      15'b001_100111011110 : VALUE=19'b0000000_110010010101;
      15'b001_100111011111 : VALUE=19'b0000000_110010010101;
      15'b001_100111100000 : VALUE=19'b0000000_110010010101;
      15'b001_100111100001 : VALUE=19'b0000000_110010010101;
      15'b001_100111100010 : VALUE=19'b0000000_110010010100;
      15'b001_100111100011 : VALUE=19'b0000000_110010010100;
      15'b001_100111100100 : VALUE=19'b0000000_110010010100;
      15'b001_100111100101 : VALUE=19'b0000000_110010010100;
      15'b001_100111100110 : VALUE=19'b0000000_110010010011;
      15'b001_100111100111 : VALUE=19'b0000000_110010010011;
      15'b001_100111101000 : VALUE=19'b0000000_110010010011;
      15'b001_100111101001 : VALUE=19'b0000000_110010010011;
      15'b001_100111101010 : VALUE=19'b0000000_110010010010;
      15'b001_100111101011 : VALUE=19'b0000000_110010010010;
      15'b001_100111101100 : VALUE=19'b0000000_110010010010;
      15'b001_100111101101 : VALUE=19'b0000000_110010010010;
      15'b001_100111101110 : VALUE=19'b0000000_110010010010;
      15'b001_100111101111 : VALUE=19'b0000000_110010010001;
      15'b001_100111110000 : VALUE=19'b0000000_110010010001;
      15'b001_100111110001 : VALUE=19'b0000000_110010010001;
      15'b001_100111110010 : VALUE=19'b0000000_110010010001;
      15'b001_100111110011 : VALUE=19'b0000000_110010010000;
      15'b001_100111110100 : VALUE=19'b0000000_110010010000;
      15'b001_100111110101 : VALUE=19'b0000000_110010010000;
      15'b001_100111110110 : VALUE=19'b0000000_110010010000;
      15'b001_100111110111 : VALUE=19'b0000000_110010001111;
      15'b001_100111111000 : VALUE=19'b0000000_110010001111;
      15'b001_100111111001 : VALUE=19'b0000000_110010001111;
      15'b001_100111111010 : VALUE=19'b0000000_110010001111;
      15'b001_100111111011 : VALUE=19'b0000000_110010001110;
      15'b001_100111111100 : VALUE=19'b0000000_110010001110;
      15'b001_100111111101 : VALUE=19'b0000000_110010001110;
      15'b001_100111111110 : VALUE=19'b0000000_110010001110;
      15'b001_100111111111 : VALUE=19'b0000000_110010001101;
      15'b001_101000000000 : VALUE=19'b0000000_110010001101;
      15'b001_101000000001 : VALUE=19'b0000000_110010001101;
      15'b001_101000000010 : VALUE=19'b0000000_110010001101;
      15'b001_101000000011 : VALUE=19'b0000000_110010001100;
      15'b001_101000000100 : VALUE=19'b0000000_110010001100;
      15'b001_101000000101 : VALUE=19'b0000000_110010001100;
      15'b001_101000000110 : VALUE=19'b0000000_110010001100;
      15'b001_101000000111 : VALUE=19'b0000000_110010001011;
      15'b001_101000001000 : VALUE=19'b0000000_110010001011;
      15'b001_101000001001 : VALUE=19'b0000000_110010001011;
      15'b001_101000001010 : VALUE=19'b0000000_110010001011;
      15'b001_101000001011 : VALUE=19'b0000000_110010001011;
      15'b001_101000001100 : VALUE=19'b0000000_110010001010;
      15'b001_101000001101 : VALUE=19'b0000000_110010001010;
      15'b001_101000001110 : VALUE=19'b0000000_110010001010;
      15'b001_101000001111 : VALUE=19'b0000000_110010001010;
      15'b001_101000010000 : VALUE=19'b0000000_110010001001;
      15'b001_101000010001 : VALUE=19'b0000000_110010001001;
      15'b001_101000010010 : VALUE=19'b0000000_110010001001;
      15'b001_101000010011 : VALUE=19'b0000000_110010001001;
      15'b001_101000010100 : VALUE=19'b0000000_110010001000;
      15'b001_101000010101 : VALUE=19'b0000000_110010001000;
      15'b001_101000010110 : VALUE=19'b0000000_110010001000;
      15'b001_101000010111 : VALUE=19'b0000000_110010001000;
      15'b001_101000011000 : VALUE=19'b0000000_110010000111;
      15'b001_101000011001 : VALUE=19'b0000000_110010000111;
      15'b001_101000011010 : VALUE=19'b0000000_110010000111;
      15'b001_101000011011 : VALUE=19'b0000000_110010000111;
      15'b001_101000011100 : VALUE=19'b0000000_110010000110;
      15'b001_101000011101 : VALUE=19'b0000000_110010000110;
      15'b001_101000011110 : VALUE=19'b0000000_110010000110;
      15'b001_101000011111 : VALUE=19'b0000000_110010000110;
      15'b001_101000100000 : VALUE=19'b0000000_110010000101;
      15'b001_101000100001 : VALUE=19'b0000000_110010000101;
      15'b001_101000100010 : VALUE=19'b0000000_110010000101;
      15'b001_101000100011 : VALUE=19'b0000000_110010000101;
      15'b001_101000100100 : VALUE=19'b0000000_110010000101;
      15'b001_101000100101 : VALUE=19'b0000000_110010000100;
      15'b001_101000100110 : VALUE=19'b0000000_110010000100;
      15'b001_101000100111 : VALUE=19'b0000000_110010000100;
      15'b001_101000101000 : VALUE=19'b0000000_110010000100;
      15'b001_101000101001 : VALUE=19'b0000000_110010000011;
      15'b001_101000101010 : VALUE=19'b0000000_110010000011;
      15'b001_101000101011 : VALUE=19'b0000000_110010000011;
      15'b001_101000101100 : VALUE=19'b0000000_110010000011;
      15'b001_101000101101 : VALUE=19'b0000000_110010000010;
      15'b001_101000101110 : VALUE=19'b0000000_110010000010;
      15'b001_101000101111 : VALUE=19'b0000000_110010000010;
      15'b001_101000110000 : VALUE=19'b0000000_110010000010;
      15'b001_101000110001 : VALUE=19'b0000000_110010000001;
      15'b001_101000110010 : VALUE=19'b0000000_110010000001;
      15'b001_101000110011 : VALUE=19'b0000000_110010000001;
      15'b001_101000110100 : VALUE=19'b0000000_110010000001;
      15'b001_101000110101 : VALUE=19'b0000000_110010000000;
      15'b001_101000110110 : VALUE=19'b0000000_110010000000;
      15'b001_101000110111 : VALUE=19'b0000000_110010000000;
      15'b001_101000111000 : VALUE=19'b0000000_110010000000;
      15'b001_101000111001 : VALUE=19'b0000000_110001111111;
      15'b001_101000111010 : VALUE=19'b0000000_110001111111;
      15'b001_101000111011 : VALUE=19'b0000000_110001111111;
      15'b001_101000111100 : VALUE=19'b0000000_110001111111;
      15'b001_101000111101 : VALUE=19'b0000000_110001111111;
      15'b001_101000111110 : VALUE=19'b0000000_110001111110;
      15'b001_101000111111 : VALUE=19'b0000000_110001111110;
      15'b001_101001000000 : VALUE=19'b0000000_110001111110;
      15'b001_101001000001 : VALUE=19'b0000000_110001111110;
      15'b001_101001000010 : VALUE=19'b0000000_110001111101;
      15'b001_101001000011 : VALUE=19'b0000000_110001111101;
      15'b001_101001000100 : VALUE=19'b0000000_110001111101;
      15'b001_101001000101 : VALUE=19'b0000000_110001111101;
      15'b001_101001000110 : VALUE=19'b0000000_110001111100;
      15'b001_101001000111 : VALUE=19'b0000000_110001111100;
      15'b001_101001001000 : VALUE=19'b0000000_110001111100;
      15'b001_101001001001 : VALUE=19'b0000000_110001111100;
      15'b001_101001001010 : VALUE=19'b0000000_110001111011;
      15'b001_101001001011 : VALUE=19'b0000000_110001111011;
      15'b001_101001001100 : VALUE=19'b0000000_110001111011;
      15'b001_101001001101 : VALUE=19'b0000000_110001111011;
      15'b001_101001001110 : VALUE=19'b0000000_110001111011;
      15'b001_101001001111 : VALUE=19'b0000000_110001111010;
      15'b001_101001010000 : VALUE=19'b0000000_110001111010;
      15'b001_101001010001 : VALUE=19'b0000000_110001111010;
      15'b001_101001010010 : VALUE=19'b0000000_110001111010;
      15'b001_101001010011 : VALUE=19'b0000000_110001111001;
      15'b001_101001010100 : VALUE=19'b0000000_110001111001;
      15'b001_101001010101 : VALUE=19'b0000000_110001111001;
      15'b001_101001010110 : VALUE=19'b0000000_110001111001;
      15'b001_101001010111 : VALUE=19'b0000000_110001111000;
      15'b001_101001011000 : VALUE=19'b0000000_110001111000;
      15'b001_101001011001 : VALUE=19'b0000000_110001111000;
      15'b001_101001011010 : VALUE=19'b0000000_110001111000;
      15'b001_101001011011 : VALUE=19'b0000000_110001110111;
      15'b001_101001011100 : VALUE=19'b0000000_110001110111;
      15'b001_101001011101 : VALUE=19'b0000000_110001110111;
      15'b001_101001011110 : VALUE=19'b0000000_110001110111;
      15'b001_101001011111 : VALUE=19'b0000000_110001110110;
      15'b001_101001100000 : VALUE=19'b0000000_110001110110;
      15'b001_101001100001 : VALUE=19'b0000000_110001110110;
      15'b001_101001100010 : VALUE=19'b0000000_110001110110;
      15'b001_101001100011 : VALUE=19'b0000000_110001110110;
      15'b001_101001100100 : VALUE=19'b0000000_110001110101;
      15'b001_101001100101 : VALUE=19'b0000000_110001110101;
      15'b001_101001100110 : VALUE=19'b0000000_110001110101;
      15'b001_101001100111 : VALUE=19'b0000000_110001110101;
      15'b001_101001101000 : VALUE=19'b0000000_110001110100;
      15'b001_101001101001 : VALUE=19'b0000000_110001110100;
      15'b001_101001101010 : VALUE=19'b0000000_110001110100;
      15'b001_101001101011 : VALUE=19'b0000000_110001110100;
      15'b001_101001101100 : VALUE=19'b0000000_110001110011;
      15'b001_101001101101 : VALUE=19'b0000000_110001110011;
      15'b001_101001101110 : VALUE=19'b0000000_110001110011;
      15'b001_101001101111 : VALUE=19'b0000000_110001110011;
      15'b001_101001110000 : VALUE=19'b0000000_110001110010;
      15'b001_101001110001 : VALUE=19'b0000000_110001110010;
      15'b001_101001110010 : VALUE=19'b0000000_110001110010;
      15'b001_101001110011 : VALUE=19'b0000000_110001110010;
      15'b001_101001110100 : VALUE=19'b0000000_110001110010;
      15'b001_101001110101 : VALUE=19'b0000000_110001110001;
      15'b001_101001110110 : VALUE=19'b0000000_110001110001;
      15'b001_101001110111 : VALUE=19'b0000000_110001110001;
      15'b001_101001111000 : VALUE=19'b0000000_110001110001;
      15'b001_101001111001 : VALUE=19'b0000000_110001110000;
      15'b001_101001111010 : VALUE=19'b0000000_110001110000;
      15'b001_101001111011 : VALUE=19'b0000000_110001110000;
      15'b001_101001111100 : VALUE=19'b0000000_110001110000;
      15'b001_101001111101 : VALUE=19'b0000000_110001101111;
      15'b001_101001111110 : VALUE=19'b0000000_110001101111;
      15'b001_101001111111 : VALUE=19'b0000000_110001101111;
      15'b001_101010000000 : VALUE=19'b0000000_110001101111;
      15'b001_101010000001 : VALUE=19'b0000000_110001101110;
      15'b001_101010000010 : VALUE=19'b0000000_110001101110;
      15'b001_101010000011 : VALUE=19'b0000000_110001101110;
      15'b001_101010000100 : VALUE=19'b0000000_110001101110;
      15'b001_101010000101 : VALUE=19'b0000000_110001101110;
      15'b001_101010000110 : VALUE=19'b0000000_110001101101;
      15'b001_101010000111 : VALUE=19'b0000000_110001101101;
      15'b001_101010001000 : VALUE=19'b0000000_110001101101;
      15'b001_101010001001 : VALUE=19'b0000000_110001101101;
      15'b001_101010001010 : VALUE=19'b0000000_110001101100;
      15'b001_101010001011 : VALUE=19'b0000000_110001101100;
      15'b001_101010001100 : VALUE=19'b0000000_110001101100;
      15'b001_101010001101 : VALUE=19'b0000000_110001101100;
      15'b001_101010001110 : VALUE=19'b0000000_110001101011;
      15'b001_101010001111 : VALUE=19'b0000000_110001101011;
      15'b001_101010010000 : VALUE=19'b0000000_110001101011;
      15'b001_101010010001 : VALUE=19'b0000000_110001101011;
      15'b001_101010010010 : VALUE=19'b0000000_110001101010;
      15'b001_101010010011 : VALUE=19'b0000000_110001101010;
      15'b001_101010010100 : VALUE=19'b0000000_110001101010;
      15'b001_101010010101 : VALUE=19'b0000000_110001101010;
      15'b001_101010010110 : VALUE=19'b0000000_110001101010;
      15'b001_101010010111 : VALUE=19'b0000000_110001101001;
      15'b001_101010011000 : VALUE=19'b0000000_110001101001;
      15'b001_101010011001 : VALUE=19'b0000000_110001101001;
      15'b001_101010011010 : VALUE=19'b0000000_110001101001;
      15'b001_101010011011 : VALUE=19'b0000000_110001101000;
      15'b001_101010011100 : VALUE=19'b0000000_110001101000;
      15'b001_101010011101 : VALUE=19'b0000000_110001101000;
      15'b001_101010011110 : VALUE=19'b0000000_110001101000;
      15'b001_101010011111 : VALUE=19'b0000000_110001100111;
      15'b001_101010100000 : VALUE=19'b0000000_110001100111;
      15'b001_101010100001 : VALUE=19'b0000000_110001100111;
      15'b001_101010100010 : VALUE=19'b0000000_110001100111;
      15'b001_101010100011 : VALUE=19'b0000000_110001100111;
      15'b001_101010100100 : VALUE=19'b0000000_110001100110;
      15'b001_101010100101 : VALUE=19'b0000000_110001100110;
      15'b001_101010100110 : VALUE=19'b0000000_110001100110;
      15'b001_101010100111 : VALUE=19'b0000000_110001100110;
      15'b001_101010101000 : VALUE=19'b0000000_110001100101;
      15'b001_101010101001 : VALUE=19'b0000000_110001100101;
      15'b001_101010101010 : VALUE=19'b0000000_110001100101;
      15'b001_101010101011 : VALUE=19'b0000000_110001100101;
      15'b001_101010101100 : VALUE=19'b0000000_110001100100;
      15'b001_101010101101 : VALUE=19'b0000000_110001100100;
      15'b001_101010101110 : VALUE=19'b0000000_110001100100;
      15'b001_101010101111 : VALUE=19'b0000000_110001100100;
      15'b001_101010110000 : VALUE=19'b0000000_110001100100;
      15'b001_101010110001 : VALUE=19'b0000000_110001100011;
      15'b001_101010110010 : VALUE=19'b0000000_110001100011;
      15'b001_101010110011 : VALUE=19'b0000000_110001100011;
      15'b001_101010110100 : VALUE=19'b0000000_110001100011;
      15'b001_101010110101 : VALUE=19'b0000000_110001100010;
      15'b001_101010110110 : VALUE=19'b0000000_110001100010;
      15'b001_101010110111 : VALUE=19'b0000000_110001100010;
      15'b001_101010111000 : VALUE=19'b0000000_110001100010;
      15'b001_101010111001 : VALUE=19'b0000000_110001100001;
      15'b001_101010111010 : VALUE=19'b0000000_110001100001;
      15'b001_101010111011 : VALUE=19'b0000000_110001100001;
      15'b001_101010111100 : VALUE=19'b0000000_110001100001;
      15'b001_101010111101 : VALUE=19'b0000000_110001100000;
      15'b001_101010111110 : VALUE=19'b0000000_110001100000;
      15'b001_101010111111 : VALUE=19'b0000000_110001100000;
      15'b001_101011000000 : VALUE=19'b0000000_110001100000;
      15'b001_101011000001 : VALUE=19'b0000000_110001100000;
      15'b001_101011000010 : VALUE=19'b0000000_110001011111;
      15'b001_101011000011 : VALUE=19'b0000000_110001011111;
      15'b001_101011000100 : VALUE=19'b0000000_110001011111;
      15'b001_101011000101 : VALUE=19'b0000000_110001011111;
      15'b001_101011000110 : VALUE=19'b0000000_110001011110;
      15'b001_101011000111 : VALUE=19'b0000000_110001011110;
      15'b001_101011001000 : VALUE=19'b0000000_110001011110;
      15'b001_101011001001 : VALUE=19'b0000000_110001011110;
      15'b001_101011001010 : VALUE=19'b0000000_110001011101;
      15'b001_101011001011 : VALUE=19'b0000000_110001011101;
      15'b001_101011001100 : VALUE=19'b0000000_110001011101;
      15'b001_101011001101 : VALUE=19'b0000000_110001011101;
      15'b001_101011001110 : VALUE=19'b0000000_110001011101;
      15'b001_101011001111 : VALUE=19'b0000000_110001011100;
      15'b001_101011010000 : VALUE=19'b0000000_110001011100;
      15'b001_101011010001 : VALUE=19'b0000000_110001011100;
      15'b001_101011010010 : VALUE=19'b0000000_110001011100;
      15'b001_101011010011 : VALUE=19'b0000000_110001011011;
      15'b001_101011010100 : VALUE=19'b0000000_110001011011;
      15'b001_101011010101 : VALUE=19'b0000000_110001011011;
      15'b001_101011010110 : VALUE=19'b0000000_110001011011;
      15'b001_101011010111 : VALUE=19'b0000000_110001011010;
      15'b001_101011011000 : VALUE=19'b0000000_110001011010;
      15'b001_101011011001 : VALUE=19'b0000000_110001011010;
      15'b001_101011011010 : VALUE=19'b0000000_110001011010;
      15'b001_101011011011 : VALUE=19'b0000000_110001011010;
      15'b001_101011011100 : VALUE=19'b0000000_110001011001;
      15'b001_101011011101 : VALUE=19'b0000000_110001011001;
      15'b001_101011011110 : VALUE=19'b0000000_110001011001;
      15'b001_101011011111 : VALUE=19'b0000000_110001011001;
      15'b001_101011100000 : VALUE=19'b0000000_110001011000;
      15'b001_101011100001 : VALUE=19'b0000000_110001011000;
      15'b001_101011100010 : VALUE=19'b0000000_110001011000;
      15'b001_101011100011 : VALUE=19'b0000000_110001011000;
      15'b001_101011100100 : VALUE=19'b0000000_110001011000;
      15'b001_101011100101 : VALUE=19'b0000000_110001010111;
      15'b001_101011100110 : VALUE=19'b0000000_110001010111;
      15'b001_101011100111 : VALUE=19'b0000000_110001010111;
      15'b001_101011101000 : VALUE=19'b0000000_110001010111;
      15'b001_101011101001 : VALUE=19'b0000000_110001010110;
      15'b001_101011101010 : VALUE=19'b0000000_110001010110;
      15'b001_101011101011 : VALUE=19'b0000000_110001010110;
      15'b001_101011101100 : VALUE=19'b0000000_110001010110;
      15'b001_101011101101 : VALUE=19'b0000000_110001010101;
      15'b001_101011101110 : VALUE=19'b0000000_110001010101;
      15'b001_101011101111 : VALUE=19'b0000000_110001010101;
      15'b001_101011110000 : VALUE=19'b0000000_110001010101;
      15'b001_101011110001 : VALUE=19'b0000000_110001010101;
      15'b001_101011110010 : VALUE=19'b0000000_110001010100;
      15'b001_101011110011 : VALUE=19'b0000000_110001010100;
      15'b001_101011110100 : VALUE=19'b0000000_110001010100;
      15'b001_101011110101 : VALUE=19'b0000000_110001010100;
      15'b001_101011110110 : VALUE=19'b0000000_110001010011;
      15'b001_101011110111 : VALUE=19'b0000000_110001010011;
      15'b001_101011111000 : VALUE=19'b0000000_110001010011;
      15'b001_101011111001 : VALUE=19'b0000000_110001010011;
      15'b001_101011111010 : VALUE=19'b0000000_110001010010;
      15'b001_101011111011 : VALUE=19'b0000000_110001010010;
      15'b001_101011111100 : VALUE=19'b0000000_110001010010;
      15'b001_101011111101 : VALUE=19'b0000000_110001010010;
      15'b001_101011111110 : VALUE=19'b0000000_110001010010;
      15'b001_101011111111 : VALUE=19'b0000000_110001010001;
      15'b001_101100000000 : VALUE=19'b0000000_110001010001;
      15'b001_101100000001 : VALUE=19'b0000000_110001010001;
      15'b001_101100000010 : VALUE=19'b0000000_110001010001;
      15'b001_101100000011 : VALUE=19'b0000000_110001010000;
      15'b001_101100000100 : VALUE=19'b0000000_110001010000;
      15'b001_101100000101 : VALUE=19'b0000000_110001010000;
      15'b001_101100000110 : VALUE=19'b0000000_110001010000;
      15'b001_101100000111 : VALUE=19'b0000000_110001010000;
      15'b001_101100001000 : VALUE=19'b0000000_110001001111;
      15'b001_101100001001 : VALUE=19'b0000000_110001001111;
      15'b001_101100001010 : VALUE=19'b0000000_110001001111;
      15'b001_101100001011 : VALUE=19'b0000000_110001001111;
      15'b001_101100001100 : VALUE=19'b0000000_110001001110;
      15'b001_101100001101 : VALUE=19'b0000000_110001001110;
      15'b001_101100001110 : VALUE=19'b0000000_110001001110;
      15'b001_101100001111 : VALUE=19'b0000000_110001001110;
      15'b001_101100010000 : VALUE=19'b0000000_110001001101;
      15'b001_101100010001 : VALUE=19'b0000000_110001001101;
      15'b001_101100010010 : VALUE=19'b0000000_110001001101;
      15'b001_101100010011 : VALUE=19'b0000000_110001001101;
      15'b001_101100010100 : VALUE=19'b0000000_110001001101;
      15'b001_101100010101 : VALUE=19'b0000000_110001001100;
      15'b001_101100010110 : VALUE=19'b0000000_110001001100;
      15'b001_101100010111 : VALUE=19'b0000000_110001001100;
      15'b001_101100011000 : VALUE=19'b0000000_110001001100;
      15'b001_101100011001 : VALUE=19'b0000000_110001001011;
      15'b001_101100011010 : VALUE=19'b0000000_110001001011;
      15'b001_101100011011 : VALUE=19'b0000000_110001001011;
      15'b001_101100011100 : VALUE=19'b0000000_110001001011;
      15'b001_101100011101 : VALUE=19'b0000000_110001001011;
      15'b001_101100011110 : VALUE=19'b0000000_110001001010;
      15'b001_101100011111 : VALUE=19'b0000000_110001001010;
      15'b001_101100100000 : VALUE=19'b0000000_110001001010;
      15'b001_101100100001 : VALUE=19'b0000000_110001001010;
      15'b001_101100100010 : VALUE=19'b0000000_110001001001;
      15'b001_101100100011 : VALUE=19'b0000000_110001001001;
      15'b001_101100100100 : VALUE=19'b0000000_110001001001;
      15'b001_101100100101 : VALUE=19'b0000000_110001001001;
      15'b001_101100100110 : VALUE=19'b0000000_110001001000;
      15'b001_101100100111 : VALUE=19'b0000000_110001001000;
      15'b001_101100101000 : VALUE=19'b0000000_110001001000;
      15'b001_101100101001 : VALUE=19'b0000000_110001001000;
      15'b001_101100101010 : VALUE=19'b0000000_110001001000;
      15'b001_101100101011 : VALUE=19'b0000000_110001000111;
      15'b001_101100101100 : VALUE=19'b0000000_110001000111;
      15'b001_101100101101 : VALUE=19'b0000000_110001000111;
      15'b001_101100101110 : VALUE=19'b0000000_110001000111;
      15'b001_101100101111 : VALUE=19'b0000000_110001000110;
      15'b001_101100110000 : VALUE=19'b0000000_110001000110;
      15'b001_101100110001 : VALUE=19'b0000000_110001000110;
      15'b001_101100110010 : VALUE=19'b0000000_110001000110;
      15'b001_101100110011 : VALUE=19'b0000000_110001000110;
      15'b001_101100110100 : VALUE=19'b0000000_110001000101;
      15'b001_101100110101 : VALUE=19'b0000000_110001000101;
      15'b001_101100110110 : VALUE=19'b0000000_110001000101;
      15'b001_101100110111 : VALUE=19'b0000000_110001000101;
      15'b001_101100111000 : VALUE=19'b0000000_110001000100;
      15'b001_101100111001 : VALUE=19'b0000000_110001000100;
      15'b001_101100111010 : VALUE=19'b0000000_110001000100;
      15'b001_101100111011 : VALUE=19'b0000000_110001000100;
      15'b001_101100111100 : VALUE=19'b0000000_110001000100;
      15'b001_101100111101 : VALUE=19'b0000000_110001000011;
      15'b001_101100111110 : VALUE=19'b0000000_110001000011;
      15'b001_101100111111 : VALUE=19'b0000000_110001000011;
      15'b001_101101000000 : VALUE=19'b0000000_110001000011;
      15'b001_101101000001 : VALUE=19'b0000000_110001000010;
      15'b001_101101000010 : VALUE=19'b0000000_110001000010;
      15'b001_101101000011 : VALUE=19'b0000000_110001000010;
      15'b001_101101000100 : VALUE=19'b0000000_110001000010;
      15'b001_101101000101 : VALUE=19'b0000000_110001000001;
      15'b001_101101000110 : VALUE=19'b0000000_110001000001;
      15'b001_101101000111 : VALUE=19'b0000000_110001000001;
      15'b001_101101001000 : VALUE=19'b0000000_110001000001;
      15'b001_101101001001 : VALUE=19'b0000000_110001000001;
      15'b001_101101001010 : VALUE=19'b0000000_110001000000;
      15'b001_101101001011 : VALUE=19'b0000000_110001000000;
      15'b001_101101001100 : VALUE=19'b0000000_110001000000;
      15'b001_101101001101 : VALUE=19'b0000000_110001000000;
      15'b001_101101001110 : VALUE=19'b0000000_110000111111;
      15'b001_101101001111 : VALUE=19'b0000000_110000111111;
      15'b001_101101010000 : VALUE=19'b0000000_110000111111;
      15'b001_101101010001 : VALUE=19'b0000000_110000111111;
      15'b001_101101010010 : VALUE=19'b0000000_110000111111;
      15'b001_101101010011 : VALUE=19'b0000000_110000111110;
      15'b001_101101010100 : VALUE=19'b0000000_110000111110;
      15'b001_101101010101 : VALUE=19'b0000000_110000111110;
      15'b001_101101010110 : VALUE=19'b0000000_110000111110;
      15'b001_101101010111 : VALUE=19'b0000000_110000111101;
      15'b001_101101011000 : VALUE=19'b0000000_110000111101;
      15'b001_101101011001 : VALUE=19'b0000000_110000111101;
      15'b001_101101011010 : VALUE=19'b0000000_110000111101;
      15'b001_101101011011 : VALUE=19'b0000000_110000111101;
      15'b001_101101011100 : VALUE=19'b0000000_110000111100;
      15'b001_101101011101 : VALUE=19'b0000000_110000111100;
      15'b001_101101011110 : VALUE=19'b0000000_110000111100;
      15'b001_101101011111 : VALUE=19'b0000000_110000111100;
      15'b001_101101100000 : VALUE=19'b0000000_110000111011;
      15'b001_101101100001 : VALUE=19'b0000000_110000111011;
      15'b001_101101100010 : VALUE=19'b0000000_110000111011;
      15'b001_101101100011 : VALUE=19'b0000000_110000111011;
      15'b001_101101100100 : VALUE=19'b0000000_110000111011;
      15'b001_101101100101 : VALUE=19'b0000000_110000111010;
      15'b001_101101100110 : VALUE=19'b0000000_110000111010;
      15'b001_101101100111 : VALUE=19'b0000000_110000111010;
      15'b001_101101101000 : VALUE=19'b0000000_110000111010;
      15'b001_101101101001 : VALUE=19'b0000000_110000111001;
      15'b001_101101101010 : VALUE=19'b0000000_110000111001;
      15'b001_101101101011 : VALUE=19'b0000000_110000111001;
      15'b001_101101101100 : VALUE=19'b0000000_110000111001;
      15'b001_101101101101 : VALUE=19'b0000000_110000111001;
      15'b001_101101101110 : VALUE=19'b0000000_110000111000;
      15'b001_101101101111 : VALUE=19'b0000000_110000111000;
      15'b001_101101110000 : VALUE=19'b0000000_110000111000;
      15'b001_101101110001 : VALUE=19'b0000000_110000111000;
      15'b001_101101110010 : VALUE=19'b0000000_110000110111;
      15'b001_101101110011 : VALUE=19'b0000000_110000110111;
      15'b001_101101110100 : VALUE=19'b0000000_110000110111;
      15'b001_101101110101 : VALUE=19'b0000000_110000110111;
      15'b001_101101110110 : VALUE=19'b0000000_110000110111;
      15'b001_101101110111 : VALUE=19'b0000000_110000110110;
      15'b001_101101111000 : VALUE=19'b0000000_110000110110;
      15'b001_101101111001 : VALUE=19'b0000000_110000110110;
      15'b001_101101111010 : VALUE=19'b0000000_110000110110;
      15'b001_101101111011 : VALUE=19'b0000000_110000110101;
      15'b001_101101111100 : VALUE=19'b0000000_110000110101;
      15'b001_101101111101 : VALUE=19'b0000000_110000110101;
      15'b001_101101111110 : VALUE=19'b0000000_110000110101;
      15'b001_101101111111 : VALUE=19'b0000000_110000110101;
      15'b001_101110000000 : VALUE=19'b0000000_110000110100;
      15'b001_101110000001 : VALUE=19'b0000000_110000110100;
      15'b001_101110000010 : VALUE=19'b0000000_110000110100;
      15'b001_101110000011 : VALUE=19'b0000000_110000110100;
      15'b001_101110000100 : VALUE=19'b0000000_110000110011;
      15'b001_101110000101 : VALUE=19'b0000000_110000110011;
      15'b001_101110000110 : VALUE=19'b0000000_110000110011;
      15'b001_101110000111 : VALUE=19'b0000000_110000110011;
      15'b001_101110001000 : VALUE=19'b0000000_110000110011;
      15'b001_101110001001 : VALUE=19'b0000000_110000110010;
      15'b001_101110001010 : VALUE=19'b0000000_110000110010;
      15'b001_101110001011 : VALUE=19'b0000000_110000110010;
      15'b001_101110001100 : VALUE=19'b0000000_110000110010;
      15'b001_101110001101 : VALUE=19'b0000000_110000110001;
      15'b001_101110001110 : VALUE=19'b0000000_110000110001;
      15'b001_101110001111 : VALUE=19'b0000000_110000110001;
      15'b001_101110010000 : VALUE=19'b0000000_110000110001;
      15'b001_101110010001 : VALUE=19'b0000000_110000110001;
      15'b001_101110010010 : VALUE=19'b0000000_110000110000;
      15'b001_101110010011 : VALUE=19'b0000000_110000110000;
      15'b001_101110010100 : VALUE=19'b0000000_110000110000;
      15'b001_101110010101 : VALUE=19'b0000000_110000110000;
      15'b001_101110010110 : VALUE=19'b0000000_110000101111;
      15'b001_101110010111 : VALUE=19'b0000000_110000101111;
      15'b001_101110011000 : VALUE=19'b0000000_110000101111;
      15'b001_101110011001 : VALUE=19'b0000000_110000101111;
      15'b001_101110011010 : VALUE=19'b0000000_110000101111;
      15'b001_101110011011 : VALUE=19'b0000000_110000101110;
      15'b001_101110011100 : VALUE=19'b0000000_110000101110;
      15'b001_101110011101 : VALUE=19'b0000000_110000101110;
      15'b001_101110011110 : VALUE=19'b0000000_110000101110;
      15'b001_101110011111 : VALUE=19'b0000000_110000101101;
      15'b001_101110100000 : VALUE=19'b0000000_110000101101;
      15'b001_101110100001 : VALUE=19'b0000000_110000101101;
      15'b001_101110100010 : VALUE=19'b0000000_110000101101;
      15'b001_101110100011 : VALUE=19'b0000000_110000101101;
      15'b001_101110100100 : VALUE=19'b0000000_110000101100;
      15'b001_101110100101 : VALUE=19'b0000000_110000101100;
      15'b001_101110100110 : VALUE=19'b0000000_110000101100;
      15'b001_101110100111 : VALUE=19'b0000000_110000101100;
      15'b001_101110101000 : VALUE=19'b0000000_110000101011;
      15'b001_101110101001 : VALUE=19'b0000000_110000101011;
      15'b001_101110101010 : VALUE=19'b0000000_110000101011;
      15'b001_101110101011 : VALUE=19'b0000000_110000101011;
      15'b001_101110101100 : VALUE=19'b0000000_110000101011;
      15'b001_101110101101 : VALUE=19'b0000000_110000101010;
      15'b001_101110101110 : VALUE=19'b0000000_110000101010;
      15'b001_101110101111 : VALUE=19'b0000000_110000101010;
      15'b001_101110110000 : VALUE=19'b0000000_110000101010;
      15'b001_101110110001 : VALUE=19'b0000000_110000101001;
      15'b001_101110110010 : VALUE=19'b0000000_110000101001;
      15'b001_101110110011 : VALUE=19'b0000000_110000101001;
      15'b001_101110110100 : VALUE=19'b0000000_110000101001;
      15'b001_101110110101 : VALUE=19'b0000000_110000101001;
      15'b001_101110110110 : VALUE=19'b0000000_110000101000;
      15'b001_101110110111 : VALUE=19'b0000000_110000101000;
      15'b001_101110111000 : VALUE=19'b0000000_110000101000;
      15'b001_101110111001 : VALUE=19'b0000000_110000101000;
      15'b001_101110111010 : VALUE=19'b0000000_110000101000;
      15'b001_101110111011 : VALUE=19'b0000000_110000100111;
      15'b001_101110111100 : VALUE=19'b0000000_110000100111;
      15'b001_101110111101 : VALUE=19'b0000000_110000100111;
      15'b001_101110111110 : VALUE=19'b0000000_110000100111;
      15'b001_101110111111 : VALUE=19'b0000000_110000100110;
      15'b001_101111000000 : VALUE=19'b0000000_110000100110;
      15'b001_101111000001 : VALUE=19'b0000000_110000100110;
      15'b001_101111000010 : VALUE=19'b0000000_110000100110;
      15'b001_101111000011 : VALUE=19'b0000000_110000100110;
      15'b001_101111000100 : VALUE=19'b0000000_110000100101;
      15'b001_101111000101 : VALUE=19'b0000000_110000100101;
      15'b001_101111000110 : VALUE=19'b0000000_110000100101;
      15'b001_101111000111 : VALUE=19'b0000000_110000100101;
      15'b001_101111001000 : VALUE=19'b0000000_110000100100;
      15'b001_101111001001 : VALUE=19'b0000000_110000100100;
      15'b001_101111001010 : VALUE=19'b0000000_110000100100;
      15'b001_101111001011 : VALUE=19'b0000000_110000100100;
      15'b001_101111001100 : VALUE=19'b0000000_110000100100;
      15'b001_101111001101 : VALUE=19'b0000000_110000100011;
      15'b001_101111001110 : VALUE=19'b0000000_110000100011;
      15'b001_101111001111 : VALUE=19'b0000000_110000100011;
      15'b001_101111010000 : VALUE=19'b0000000_110000100011;
      15'b001_101111010001 : VALUE=19'b0000000_110000100010;
      15'b001_101111010010 : VALUE=19'b0000000_110000100010;
      15'b001_101111010011 : VALUE=19'b0000000_110000100010;
      15'b001_101111010100 : VALUE=19'b0000000_110000100010;
      15'b001_101111010101 : VALUE=19'b0000000_110000100010;
      15'b001_101111010110 : VALUE=19'b0000000_110000100001;
      15'b001_101111010111 : VALUE=19'b0000000_110000100001;
      15'b001_101111011000 : VALUE=19'b0000000_110000100001;
      15'b001_101111011001 : VALUE=19'b0000000_110000100001;
      15'b001_101111011010 : VALUE=19'b0000000_110000100001;
      15'b001_101111011011 : VALUE=19'b0000000_110000100000;
      15'b001_101111011100 : VALUE=19'b0000000_110000100000;
      15'b001_101111011101 : VALUE=19'b0000000_110000100000;
      15'b001_101111011110 : VALUE=19'b0000000_110000100000;
      15'b001_101111011111 : VALUE=19'b0000000_110000011111;
      15'b001_101111100000 : VALUE=19'b0000000_110000011111;
      15'b001_101111100001 : VALUE=19'b0000000_110000011111;
      15'b001_101111100010 : VALUE=19'b0000000_110000011111;
      15'b001_101111100011 : VALUE=19'b0000000_110000011111;
      15'b001_101111100100 : VALUE=19'b0000000_110000011110;
      15'b001_101111100101 : VALUE=19'b0000000_110000011110;
      15'b001_101111100110 : VALUE=19'b0000000_110000011110;
      15'b001_101111100111 : VALUE=19'b0000000_110000011110;
      15'b001_101111101000 : VALUE=19'b0000000_110000011101;
      15'b001_101111101001 : VALUE=19'b0000000_110000011101;
      15'b001_101111101010 : VALUE=19'b0000000_110000011101;
      15'b001_101111101011 : VALUE=19'b0000000_110000011101;
      15'b001_101111101100 : VALUE=19'b0000000_110000011101;
      15'b001_101111101101 : VALUE=19'b0000000_110000011100;
      15'b001_101111101110 : VALUE=19'b0000000_110000011100;
      15'b001_101111101111 : VALUE=19'b0000000_110000011100;
      15'b001_101111110000 : VALUE=19'b0000000_110000011100;
      15'b001_101111110001 : VALUE=19'b0000000_110000011100;
      15'b001_101111110010 : VALUE=19'b0000000_110000011011;
      15'b001_101111110011 : VALUE=19'b0000000_110000011011;
      15'b001_101111110100 : VALUE=19'b0000000_110000011011;
      15'b001_101111110101 : VALUE=19'b0000000_110000011011;
      15'b001_101111110110 : VALUE=19'b0000000_110000011010;
      15'b001_101111110111 : VALUE=19'b0000000_110000011010;
      15'b001_101111111000 : VALUE=19'b0000000_110000011010;
      15'b001_101111111001 : VALUE=19'b0000000_110000011010;
      15'b001_101111111010 : VALUE=19'b0000000_110000011010;
      15'b001_101111111011 : VALUE=19'b0000000_110000011001;
      15'b001_101111111100 : VALUE=19'b0000000_110000011001;
      15'b001_101111111101 : VALUE=19'b0000000_110000011001;
      15'b001_101111111110 : VALUE=19'b0000000_110000011001;
      15'b001_101111111111 : VALUE=19'b0000000_110000011001;
      15'b001_110000000000 : VALUE=19'b0000000_110000011000;
      15'b001_110000000001 : VALUE=19'b0000000_110000011000;
      15'b001_110000000010 : VALUE=19'b0000000_110000011000;
      15'b001_110000000011 : VALUE=19'b0000000_110000011000;
      15'b001_110000000100 : VALUE=19'b0000000_110000010111;
      15'b001_110000000101 : VALUE=19'b0000000_110000010111;
      15'b001_110000000110 : VALUE=19'b0000000_110000010111;
      15'b001_110000000111 : VALUE=19'b0000000_110000010111;
      15'b001_110000001000 : VALUE=19'b0000000_110000010111;
      15'b001_110000001001 : VALUE=19'b0000000_110000010110;
      15'b001_110000001010 : VALUE=19'b0000000_110000010110;
      15'b001_110000001011 : VALUE=19'b0000000_110000010110;
      15'b001_110000001100 : VALUE=19'b0000000_110000010110;
      15'b001_110000001101 : VALUE=19'b0000000_110000010101;
      15'b001_110000001110 : VALUE=19'b0000000_110000010101;
      15'b001_110000001111 : VALUE=19'b0000000_110000010101;
      15'b001_110000010000 : VALUE=19'b0000000_110000010101;
      15'b001_110000010001 : VALUE=19'b0000000_110000010101;
      15'b001_110000010010 : VALUE=19'b0000000_110000010100;
      15'b001_110000010011 : VALUE=19'b0000000_110000010100;
      15'b001_110000010100 : VALUE=19'b0000000_110000010100;
      15'b001_110000010101 : VALUE=19'b0000000_110000010100;
      15'b001_110000010110 : VALUE=19'b0000000_110000010100;
      15'b001_110000010111 : VALUE=19'b0000000_110000010011;
      15'b001_110000011000 : VALUE=19'b0000000_110000010011;
      15'b001_110000011001 : VALUE=19'b0000000_110000010011;
      15'b001_110000011010 : VALUE=19'b0000000_110000010011;
      15'b001_110000011011 : VALUE=19'b0000000_110000010010;
      15'b001_110000011100 : VALUE=19'b0000000_110000010010;
      15'b001_110000011101 : VALUE=19'b0000000_110000010010;
      15'b001_110000011110 : VALUE=19'b0000000_110000010010;
      15'b001_110000011111 : VALUE=19'b0000000_110000010010;
      15'b001_110000100000 : VALUE=19'b0000000_110000010001;
      15'b001_110000100001 : VALUE=19'b0000000_110000010001;
      15'b001_110000100010 : VALUE=19'b0000000_110000010001;
      15'b001_110000100011 : VALUE=19'b0000000_110000010001;
      15'b001_110000100100 : VALUE=19'b0000000_110000010001;
      15'b001_110000100101 : VALUE=19'b0000000_110000010000;
      15'b001_110000100110 : VALUE=19'b0000000_110000010000;
      15'b001_110000100111 : VALUE=19'b0000000_110000010000;
      15'b001_110000101000 : VALUE=19'b0000000_110000010000;
      15'b001_110000101001 : VALUE=19'b0000000_110000001111;
      15'b001_110000101010 : VALUE=19'b0000000_110000001111;
      15'b001_110000101011 : VALUE=19'b0000000_110000001111;
      15'b001_110000101100 : VALUE=19'b0000000_110000001111;
      15'b001_110000101101 : VALUE=19'b0000000_110000001111;
      15'b001_110000101110 : VALUE=19'b0000000_110000001110;
      15'b001_110000101111 : VALUE=19'b0000000_110000001110;
      15'b001_110000110000 : VALUE=19'b0000000_110000001110;
      15'b001_110000110001 : VALUE=19'b0000000_110000001110;
      15'b001_110000110010 : VALUE=19'b0000000_110000001110;
      15'b001_110000110011 : VALUE=19'b0000000_110000001101;
      15'b001_110000110100 : VALUE=19'b0000000_110000001101;
      15'b001_110000110101 : VALUE=19'b0000000_110000001101;
      15'b001_110000110110 : VALUE=19'b0000000_110000001101;
      15'b001_110000110111 : VALUE=19'b0000000_110000001100;
      15'b001_110000111000 : VALUE=19'b0000000_110000001100;
      15'b001_110000111001 : VALUE=19'b0000000_110000001100;
      15'b001_110000111010 : VALUE=19'b0000000_110000001100;
      15'b001_110000111011 : VALUE=19'b0000000_110000001100;
      15'b001_110000111100 : VALUE=19'b0000000_110000001011;
      15'b001_110000111101 : VALUE=19'b0000000_110000001011;
      15'b001_110000111110 : VALUE=19'b0000000_110000001011;
      15'b001_110000111111 : VALUE=19'b0000000_110000001011;
      15'b001_110001000000 : VALUE=19'b0000000_110000001011;
      15'b001_110001000001 : VALUE=19'b0000000_110000001010;
      15'b001_110001000010 : VALUE=19'b0000000_110000001010;
      15'b001_110001000011 : VALUE=19'b0000000_110000001010;
      15'b001_110001000100 : VALUE=19'b0000000_110000001010;
      15'b001_110001000101 : VALUE=19'b0000000_110000001001;
      15'b001_110001000110 : VALUE=19'b0000000_110000001001;
      15'b001_110001000111 : VALUE=19'b0000000_110000001001;
      15'b001_110001001000 : VALUE=19'b0000000_110000001001;
      15'b001_110001001001 : VALUE=19'b0000000_110000001001;
      15'b001_110001001010 : VALUE=19'b0000000_110000001000;
      15'b001_110001001011 : VALUE=19'b0000000_110000001000;
      15'b001_110001001100 : VALUE=19'b0000000_110000001000;
      15'b001_110001001101 : VALUE=19'b0000000_110000001000;
      15'b001_110001001110 : VALUE=19'b0000000_110000001000;
      15'b001_110001001111 : VALUE=19'b0000000_110000000111;
      15'b001_110001010000 : VALUE=19'b0000000_110000000111;
      15'b001_110001010001 : VALUE=19'b0000000_110000000111;
      15'b001_110001010010 : VALUE=19'b0000000_110000000111;
      15'b001_110001010011 : VALUE=19'b0000000_110000000111;
      15'b001_110001010100 : VALUE=19'b0000000_110000000110;
      15'b001_110001010101 : VALUE=19'b0000000_110000000110;
      15'b001_110001010110 : VALUE=19'b0000000_110000000110;
      15'b001_110001010111 : VALUE=19'b0000000_110000000110;
      15'b001_110001011000 : VALUE=19'b0000000_110000000101;
      15'b001_110001011001 : VALUE=19'b0000000_110000000101;
      15'b001_110001011010 : VALUE=19'b0000000_110000000101;
      15'b001_110001011011 : VALUE=19'b0000000_110000000101;
      15'b001_110001011100 : VALUE=19'b0000000_110000000101;
      15'b001_110001011101 : VALUE=19'b0000000_110000000100;
      15'b001_110001011110 : VALUE=19'b0000000_110000000100;
      15'b001_110001011111 : VALUE=19'b0000000_110000000100;
      15'b001_110001100000 : VALUE=19'b0000000_110000000100;
      15'b001_110001100001 : VALUE=19'b0000000_110000000100;
      15'b001_110001100010 : VALUE=19'b0000000_110000000011;
      15'b001_110001100011 : VALUE=19'b0000000_110000000011;
      15'b001_110001100100 : VALUE=19'b0000000_110000000011;
      15'b001_110001100101 : VALUE=19'b0000000_110000000011;
      15'b001_110001100110 : VALUE=19'b0000000_110000000010;
      15'b001_110001100111 : VALUE=19'b0000000_110000000010;
      15'b001_110001101000 : VALUE=19'b0000000_110000000010;
      15'b001_110001101001 : VALUE=19'b0000000_110000000010;
      15'b001_110001101010 : VALUE=19'b0000000_110000000010;
      15'b001_110001101011 : VALUE=19'b0000000_110000000001;
      15'b001_110001101100 : VALUE=19'b0000000_110000000001;
      15'b001_110001101101 : VALUE=19'b0000000_110000000001;
      15'b001_110001101110 : VALUE=19'b0000000_110000000001;
      15'b001_110001101111 : VALUE=19'b0000000_110000000001;
      15'b001_110001110000 : VALUE=19'b0000000_110000000000;
      15'b001_110001110001 : VALUE=19'b0000000_110000000000;
      15'b001_110001110010 : VALUE=19'b0000000_110000000000;
      15'b001_110001110011 : VALUE=19'b0000000_110000000000;
      15'b001_110001110100 : VALUE=19'b0000000_110000000000;
      15'b001_110001110101 : VALUE=19'b0000000_101111111111;
      15'b001_110001110110 : VALUE=19'b0000000_101111111111;
      15'b001_110001110111 : VALUE=19'b0000000_101111111111;
      15'b001_110001111000 : VALUE=19'b0000000_101111111111;
      15'b001_110001111001 : VALUE=19'b0000000_101111111110;
      15'b001_110001111010 : VALUE=19'b0000000_101111111110;
      15'b001_110001111011 : VALUE=19'b0000000_101111111110;
      15'b001_110001111100 : VALUE=19'b0000000_101111111110;
      15'b001_110001111101 : VALUE=19'b0000000_101111111110;
      15'b001_110001111110 : VALUE=19'b0000000_101111111101;
      15'b001_110001111111 : VALUE=19'b0000000_101111111101;
      15'b001_110010000000 : VALUE=19'b0000000_101111111101;
      15'b001_110010000001 : VALUE=19'b0000000_101111111101;
      15'b001_110010000010 : VALUE=19'b0000000_101111111101;
      15'b001_110010000011 : VALUE=19'b0000000_101111111100;
      15'b001_110010000100 : VALUE=19'b0000000_101111111100;
      15'b001_110010000101 : VALUE=19'b0000000_101111111100;
      15'b001_110010000110 : VALUE=19'b0000000_101111111100;
      15'b001_110010000111 : VALUE=19'b0000000_101111111100;
      15'b001_110010001000 : VALUE=19'b0000000_101111111011;
      15'b001_110010001001 : VALUE=19'b0000000_101111111011;
      15'b001_110010001010 : VALUE=19'b0000000_101111111011;
      15'b001_110010001011 : VALUE=19'b0000000_101111111011;
      15'b001_110010001100 : VALUE=19'b0000000_101111111010;
      15'b001_110010001101 : VALUE=19'b0000000_101111111010;
      15'b001_110010001110 : VALUE=19'b0000000_101111111010;
      15'b001_110010001111 : VALUE=19'b0000000_101111111010;
      15'b001_110010010000 : VALUE=19'b0000000_101111111010;
      15'b001_110010010001 : VALUE=19'b0000000_101111111001;
      15'b001_110010010010 : VALUE=19'b0000000_101111111001;
      15'b001_110010010011 : VALUE=19'b0000000_101111111001;
      15'b001_110010010100 : VALUE=19'b0000000_101111111001;
      15'b001_110010010101 : VALUE=19'b0000000_101111111001;
      15'b001_110010010110 : VALUE=19'b0000000_101111111000;
      15'b001_110010010111 : VALUE=19'b0000000_101111111000;
      15'b001_110010011000 : VALUE=19'b0000000_101111111000;
      15'b001_110010011001 : VALUE=19'b0000000_101111111000;
      15'b001_110010011010 : VALUE=19'b0000000_101111111000;
      15'b001_110010011011 : VALUE=19'b0000000_101111110111;
      15'b001_110010011100 : VALUE=19'b0000000_101111110111;
      15'b001_110010011101 : VALUE=19'b0000000_101111110111;
      15'b001_110010011110 : VALUE=19'b0000000_101111110111;
      15'b001_110010011111 : VALUE=19'b0000000_101111110111;
      15'b001_110010100000 : VALUE=19'b0000000_101111110110;
      15'b001_110010100001 : VALUE=19'b0000000_101111110110;
      15'b001_110010100010 : VALUE=19'b0000000_101111110110;
      15'b001_110010100011 : VALUE=19'b0000000_101111110110;
      15'b001_110010100100 : VALUE=19'b0000000_101111110101;
      15'b001_110010100101 : VALUE=19'b0000000_101111110101;
      15'b001_110010100110 : VALUE=19'b0000000_101111110101;
      15'b001_110010100111 : VALUE=19'b0000000_101111110101;
      15'b001_110010101000 : VALUE=19'b0000000_101111110101;
      15'b001_110010101001 : VALUE=19'b0000000_101111110100;
      15'b001_110010101010 : VALUE=19'b0000000_101111110100;
      15'b001_110010101011 : VALUE=19'b0000000_101111110100;
      15'b001_110010101100 : VALUE=19'b0000000_101111110100;
      15'b001_110010101101 : VALUE=19'b0000000_101111110100;
      15'b001_110010101110 : VALUE=19'b0000000_101111110011;
      15'b001_110010101111 : VALUE=19'b0000000_101111110011;
      15'b001_110010110000 : VALUE=19'b0000000_101111110011;
      15'b001_110010110001 : VALUE=19'b0000000_101111110011;
      15'b001_110010110010 : VALUE=19'b0000000_101111110011;
      15'b001_110010110011 : VALUE=19'b0000000_101111110010;
      15'b001_110010110100 : VALUE=19'b0000000_101111110010;
      15'b001_110010110101 : VALUE=19'b0000000_101111110010;
      15'b001_110010110110 : VALUE=19'b0000000_101111110010;
      15'b001_110010110111 : VALUE=19'b0000000_101111110010;
      15'b001_110010111000 : VALUE=19'b0000000_101111110001;
      15'b001_110010111001 : VALUE=19'b0000000_101111110001;
      15'b001_110010111010 : VALUE=19'b0000000_101111110001;
      15'b001_110010111011 : VALUE=19'b0000000_101111110001;
      15'b001_110010111100 : VALUE=19'b0000000_101111110000;
      15'b001_110010111101 : VALUE=19'b0000000_101111110000;
      15'b001_110010111110 : VALUE=19'b0000000_101111110000;
      15'b001_110010111111 : VALUE=19'b0000000_101111110000;
      15'b001_110011000000 : VALUE=19'b0000000_101111110000;
      15'b001_110011000001 : VALUE=19'b0000000_101111101111;
      15'b001_110011000010 : VALUE=19'b0000000_101111101111;
      15'b001_110011000011 : VALUE=19'b0000000_101111101111;
      15'b001_110011000100 : VALUE=19'b0000000_101111101111;
      15'b001_110011000101 : VALUE=19'b0000000_101111101111;
      15'b001_110011000110 : VALUE=19'b0000000_101111101110;
      15'b001_110011000111 : VALUE=19'b0000000_101111101110;
      15'b001_110011001000 : VALUE=19'b0000000_101111101110;
      15'b001_110011001001 : VALUE=19'b0000000_101111101110;
      15'b001_110011001010 : VALUE=19'b0000000_101111101110;
      15'b001_110011001011 : VALUE=19'b0000000_101111101101;
      15'b001_110011001100 : VALUE=19'b0000000_101111101101;
      15'b001_110011001101 : VALUE=19'b0000000_101111101101;
      15'b001_110011001110 : VALUE=19'b0000000_101111101101;
      15'b001_110011001111 : VALUE=19'b0000000_101111101101;
      15'b001_110011010000 : VALUE=19'b0000000_101111101100;
      15'b001_110011010001 : VALUE=19'b0000000_101111101100;
      15'b001_110011010010 : VALUE=19'b0000000_101111101100;
      15'b001_110011010011 : VALUE=19'b0000000_101111101100;
      15'b001_110011010100 : VALUE=19'b0000000_101111101011;
      15'b001_110011010101 : VALUE=19'b0000000_101111101011;
      15'b001_110011010110 : VALUE=19'b0000000_101111101011;
      15'b001_110011010111 : VALUE=19'b0000000_101111101011;
      15'b001_110011011000 : VALUE=19'b0000000_101111101011;
      15'b001_110011011001 : VALUE=19'b0000000_101111101010;
      15'b001_110011011010 : VALUE=19'b0000000_101111101010;
      15'b001_110011011011 : VALUE=19'b0000000_101111101010;
      15'b001_110011011100 : VALUE=19'b0000000_101111101010;
      15'b001_110011011101 : VALUE=19'b0000000_101111101010;
      15'b001_110011011110 : VALUE=19'b0000000_101111101001;
      15'b001_110011011111 : VALUE=19'b0000000_101111101001;
      15'b001_110011100000 : VALUE=19'b0000000_101111101001;
      15'b001_110011100001 : VALUE=19'b0000000_101111101001;
      15'b001_110011100010 : VALUE=19'b0000000_101111101001;
      15'b001_110011100011 : VALUE=19'b0000000_101111101000;
      15'b001_110011100100 : VALUE=19'b0000000_101111101000;
      15'b001_110011100101 : VALUE=19'b0000000_101111101000;
      15'b001_110011100110 : VALUE=19'b0000000_101111101000;
      15'b001_110011100111 : VALUE=19'b0000000_101111101000;
      15'b001_110011101000 : VALUE=19'b0000000_101111100111;
      15'b001_110011101001 : VALUE=19'b0000000_101111100111;
      15'b001_110011101010 : VALUE=19'b0000000_101111100111;
      15'b001_110011101011 : VALUE=19'b0000000_101111100111;
      15'b001_110011101100 : VALUE=19'b0000000_101111100111;
      15'b001_110011101101 : VALUE=19'b0000000_101111100110;
      15'b001_110011101110 : VALUE=19'b0000000_101111100110;
      15'b001_110011101111 : VALUE=19'b0000000_101111100110;
      15'b001_110011110000 : VALUE=19'b0000000_101111100110;
      15'b001_110011110001 : VALUE=19'b0000000_101111100110;
      15'b001_110011110010 : VALUE=19'b0000000_101111100101;
      15'b001_110011110011 : VALUE=19'b0000000_101111100101;
      15'b001_110011110100 : VALUE=19'b0000000_101111100101;
      15'b001_110011110101 : VALUE=19'b0000000_101111100101;
      15'b001_110011110110 : VALUE=19'b0000000_101111100100;
      15'b001_110011110111 : VALUE=19'b0000000_101111100100;
      15'b001_110011111000 : VALUE=19'b0000000_101111100100;
      15'b001_110011111001 : VALUE=19'b0000000_101111100100;
      15'b001_110011111010 : VALUE=19'b0000000_101111100100;
      15'b001_110011111011 : VALUE=19'b0000000_101111100011;
      15'b001_110011111100 : VALUE=19'b0000000_101111100011;
      15'b001_110011111101 : VALUE=19'b0000000_101111100011;
      15'b001_110011111110 : VALUE=19'b0000000_101111100011;
      15'b001_110011111111 : VALUE=19'b0000000_101111100011;
      15'b001_110100000000 : VALUE=19'b0000000_101111100010;
      15'b001_110100000001 : VALUE=19'b0000000_101111100010;
      15'b001_110100000010 : VALUE=19'b0000000_101111100010;
      15'b001_110100000011 : VALUE=19'b0000000_101111100010;
      15'b001_110100000100 : VALUE=19'b0000000_101111100010;
      15'b001_110100000101 : VALUE=19'b0000000_101111100001;
      15'b001_110100000110 : VALUE=19'b0000000_101111100001;
      15'b001_110100000111 : VALUE=19'b0000000_101111100001;
      15'b001_110100001000 : VALUE=19'b0000000_101111100001;
      15'b001_110100001001 : VALUE=19'b0000000_101111100001;
      15'b001_110100001010 : VALUE=19'b0000000_101111100000;
      15'b001_110100001011 : VALUE=19'b0000000_101111100000;
      15'b001_110100001100 : VALUE=19'b0000000_101111100000;
      15'b001_110100001101 : VALUE=19'b0000000_101111100000;
      15'b001_110100001110 : VALUE=19'b0000000_101111100000;
      15'b001_110100001111 : VALUE=19'b0000000_101111011111;
      15'b001_110100010000 : VALUE=19'b0000000_101111011111;
      15'b001_110100010001 : VALUE=19'b0000000_101111011111;
      15'b001_110100010010 : VALUE=19'b0000000_101111011111;
      15'b001_110100010011 : VALUE=19'b0000000_101111011111;
      15'b001_110100010100 : VALUE=19'b0000000_101111011110;
      15'b001_110100010101 : VALUE=19'b0000000_101111011110;
      15'b001_110100010110 : VALUE=19'b0000000_101111011110;
      15'b001_110100010111 : VALUE=19'b0000000_101111011110;
      15'b001_110100011000 : VALUE=19'b0000000_101111011110;
      15'b001_110100011001 : VALUE=19'b0000000_101111011101;
      15'b001_110100011010 : VALUE=19'b0000000_101111011101;
      15'b001_110100011011 : VALUE=19'b0000000_101111011101;
      15'b001_110100011100 : VALUE=19'b0000000_101111011101;
      15'b001_110100011101 : VALUE=19'b0000000_101111011101;
      15'b001_110100011110 : VALUE=19'b0000000_101111011100;
      15'b001_110100011111 : VALUE=19'b0000000_101111011100;
      15'b001_110100100000 : VALUE=19'b0000000_101111011100;
      15'b001_110100100001 : VALUE=19'b0000000_101111011100;
      15'b001_110100100010 : VALUE=19'b0000000_101111011011;
      15'b001_110100100011 : VALUE=19'b0000000_101111011011;
      15'b001_110100100100 : VALUE=19'b0000000_101111011011;
      15'b001_110100100101 : VALUE=19'b0000000_101111011011;
      15'b001_110100100110 : VALUE=19'b0000000_101111011011;
      15'b001_110100100111 : VALUE=19'b0000000_101111011010;
      15'b001_110100101000 : VALUE=19'b0000000_101111011010;
      15'b001_110100101001 : VALUE=19'b0000000_101111011010;
      15'b001_110100101010 : VALUE=19'b0000000_101111011010;
      15'b001_110100101011 : VALUE=19'b0000000_101111011010;
      15'b001_110100101100 : VALUE=19'b0000000_101111011001;
      15'b001_110100101101 : VALUE=19'b0000000_101111011001;
      15'b001_110100101110 : VALUE=19'b0000000_101111011001;
      15'b001_110100101111 : VALUE=19'b0000000_101111011001;
      15'b001_110100110000 : VALUE=19'b0000000_101111011001;
      15'b001_110100110001 : VALUE=19'b0000000_101111011000;
      15'b001_110100110010 : VALUE=19'b0000000_101111011000;
      15'b001_110100110011 : VALUE=19'b0000000_101111011000;
      15'b001_110100110100 : VALUE=19'b0000000_101111011000;
      15'b001_110100110101 : VALUE=19'b0000000_101111011000;
      15'b001_110100110110 : VALUE=19'b0000000_101111010111;
      15'b001_110100110111 : VALUE=19'b0000000_101111010111;
      15'b001_110100111000 : VALUE=19'b0000000_101111010111;
      15'b001_110100111001 : VALUE=19'b0000000_101111010111;
      15'b001_110100111010 : VALUE=19'b0000000_101111010111;
      15'b001_110100111011 : VALUE=19'b0000000_101111010110;
      15'b001_110100111100 : VALUE=19'b0000000_101111010110;
      15'b001_110100111101 : VALUE=19'b0000000_101111010110;
      15'b001_110100111110 : VALUE=19'b0000000_101111010110;
      15'b001_110100111111 : VALUE=19'b0000000_101111010110;
      15'b001_110101000000 : VALUE=19'b0000000_101111010101;
      15'b001_110101000001 : VALUE=19'b0000000_101111010101;
      15'b001_110101000010 : VALUE=19'b0000000_101111010101;
      15'b001_110101000011 : VALUE=19'b0000000_101111010101;
      15'b001_110101000100 : VALUE=19'b0000000_101111010101;
      15'b001_110101000101 : VALUE=19'b0000000_101111010100;
      15'b001_110101000110 : VALUE=19'b0000000_101111010100;
      15'b001_110101000111 : VALUE=19'b0000000_101111010100;
      15'b001_110101001000 : VALUE=19'b0000000_101111010100;
      15'b001_110101001001 : VALUE=19'b0000000_101111010100;
      15'b001_110101001010 : VALUE=19'b0000000_101111010011;
      15'b001_110101001011 : VALUE=19'b0000000_101111010011;
      15'b001_110101001100 : VALUE=19'b0000000_101111010011;
      15'b001_110101001101 : VALUE=19'b0000000_101111010011;
      15'b001_110101001110 : VALUE=19'b0000000_101111010011;
      15'b001_110101001111 : VALUE=19'b0000000_101111010010;
      15'b001_110101010000 : VALUE=19'b0000000_101111010010;
      15'b001_110101010001 : VALUE=19'b0000000_101111010010;
      15'b001_110101010010 : VALUE=19'b0000000_101111010010;
      15'b001_110101010011 : VALUE=19'b0000000_101111010010;
      15'b001_110101010100 : VALUE=19'b0000000_101111010001;
      15'b001_110101010101 : VALUE=19'b0000000_101111010001;
      15'b001_110101010110 : VALUE=19'b0000000_101111010001;
      15'b001_110101010111 : VALUE=19'b0000000_101111010001;
      15'b001_110101011000 : VALUE=19'b0000000_101111010001;
      15'b001_110101011001 : VALUE=19'b0000000_101111010000;
      15'b001_110101011010 : VALUE=19'b0000000_101111010000;
      15'b001_110101011011 : VALUE=19'b0000000_101111010000;
      15'b001_110101011100 : VALUE=19'b0000000_101111010000;
      15'b001_110101011101 : VALUE=19'b0000000_101111010000;
      15'b001_110101011110 : VALUE=19'b0000000_101111001111;
      15'b001_110101011111 : VALUE=19'b0000000_101111001111;
      15'b001_110101100000 : VALUE=19'b0000000_101111001111;
      15'b001_110101100001 : VALUE=19'b0000000_101111001111;
      15'b001_110101100010 : VALUE=19'b0000000_101111001111;
      15'b001_110101100011 : VALUE=19'b0000000_101111001110;
      15'b001_110101100100 : VALUE=19'b0000000_101111001110;
      15'b001_110101100101 : VALUE=19'b0000000_101111001110;
      15'b001_110101100110 : VALUE=19'b0000000_101111001110;
      15'b001_110101100111 : VALUE=19'b0000000_101111001110;
      15'b001_110101101000 : VALUE=19'b0000000_101111001101;
      15'b001_110101101001 : VALUE=19'b0000000_101111001101;
      15'b001_110101101010 : VALUE=19'b0000000_101111001101;
      15'b001_110101101011 : VALUE=19'b0000000_101111001101;
      15'b001_110101101100 : VALUE=19'b0000000_101111001101;
      15'b001_110101101101 : VALUE=19'b0000000_101111001100;
      15'b001_110101101110 : VALUE=19'b0000000_101111001100;
      15'b001_110101101111 : VALUE=19'b0000000_101111001100;
      15'b001_110101110000 : VALUE=19'b0000000_101111001100;
      15'b001_110101110001 : VALUE=19'b0000000_101111001100;
      15'b001_110101110010 : VALUE=19'b0000000_101111001011;
      15'b001_110101110011 : VALUE=19'b0000000_101111001011;
      15'b001_110101110100 : VALUE=19'b0000000_101111001011;
      15'b001_110101110101 : VALUE=19'b0000000_101111001011;
      15'b001_110101110110 : VALUE=19'b0000000_101111001011;
      15'b001_110101110111 : VALUE=19'b0000000_101111001010;
      15'b001_110101111000 : VALUE=19'b0000000_101111001010;
      15'b001_110101111001 : VALUE=19'b0000000_101111001010;
      15'b001_110101111010 : VALUE=19'b0000000_101111001010;
      15'b001_110101111011 : VALUE=19'b0000000_101111001010;
      15'b001_110101111100 : VALUE=19'b0000000_101111001001;
      15'b001_110101111101 : VALUE=19'b0000000_101111001001;
      15'b001_110101111110 : VALUE=19'b0000000_101111001001;
      15'b001_110101111111 : VALUE=19'b0000000_101111001001;
      15'b001_110110000000 : VALUE=19'b0000000_101111001001;
      15'b001_110110000001 : VALUE=19'b0000000_101111001000;
      15'b001_110110000010 : VALUE=19'b0000000_101111001000;
      15'b001_110110000011 : VALUE=19'b0000000_101111001000;
      15'b001_110110000100 : VALUE=19'b0000000_101111001000;
      15'b001_110110000101 : VALUE=19'b0000000_101111001000;
      15'b001_110110000110 : VALUE=19'b0000000_101111000111;
      15'b001_110110000111 : VALUE=19'b0000000_101111000111;
      15'b001_110110001000 : VALUE=19'b0000000_101111000111;
      15'b001_110110001001 : VALUE=19'b0000000_101111000111;
      15'b001_110110001010 : VALUE=19'b0000000_101111000111;
      15'b001_110110001011 : VALUE=19'b0000000_101111000110;
      15'b001_110110001100 : VALUE=19'b0000000_101111000110;
      15'b001_110110001101 : VALUE=19'b0000000_101111000110;
      15'b001_110110001110 : VALUE=19'b0000000_101111000110;
      15'b001_110110001111 : VALUE=19'b0000000_101111000110;
      15'b001_110110010000 : VALUE=19'b0000000_101111000101;
      15'b001_110110010001 : VALUE=19'b0000000_101111000101;
      15'b001_110110010010 : VALUE=19'b0000000_101111000101;
      15'b001_110110010011 : VALUE=19'b0000000_101111000101;
      15'b001_110110010100 : VALUE=19'b0000000_101111000101;
      15'b001_110110010101 : VALUE=19'b0000000_101111000100;
      15'b001_110110010110 : VALUE=19'b0000000_101111000100;
      15'b001_110110010111 : VALUE=19'b0000000_101111000100;
      15'b001_110110011000 : VALUE=19'b0000000_101111000100;
      15'b001_110110011001 : VALUE=19'b0000000_101111000100;
      15'b001_110110011010 : VALUE=19'b0000000_101111000011;
      15'b001_110110011011 : VALUE=19'b0000000_101111000011;
      15'b001_110110011100 : VALUE=19'b0000000_101111000011;
      15'b001_110110011101 : VALUE=19'b0000000_101111000011;
      15'b001_110110011110 : VALUE=19'b0000000_101111000011;
      15'b001_110110011111 : VALUE=19'b0000000_101111000010;
      15'b001_110110100000 : VALUE=19'b0000000_101111000010;
      15'b001_110110100001 : VALUE=19'b0000000_101111000010;
      15'b001_110110100010 : VALUE=19'b0000000_101111000010;
      15'b001_110110100011 : VALUE=19'b0000000_101111000010;
      15'b001_110110100100 : VALUE=19'b0000000_101111000001;
      15'b001_110110100101 : VALUE=19'b0000000_101111000001;
      15'b001_110110100110 : VALUE=19'b0000000_101111000001;
      15'b001_110110100111 : VALUE=19'b0000000_101111000001;
      15'b001_110110101000 : VALUE=19'b0000000_101111000001;
      15'b001_110110101001 : VALUE=19'b0000000_101111000000;
      15'b001_110110101010 : VALUE=19'b0000000_101111000000;
      15'b001_110110101011 : VALUE=19'b0000000_101111000000;
      15'b001_110110101100 : VALUE=19'b0000000_101111000000;
      15'b001_110110101101 : VALUE=19'b0000000_101111000000;
      15'b001_110110101110 : VALUE=19'b0000000_101110111111;
      15'b001_110110101111 : VALUE=19'b0000000_101110111111;
      15'b001_110110110000 : VALUE=19'b0000000_101110111111;
      15'b001_110110110001 : VALUE=19'b0000000_101110111111;
      15'b001_110110110010 : VALUE=19'b0000000_101110111111;
      15'b001_110110110011 : VALUE=19'b0000000_101110111110;
      15'b001_110110110100 : VALUE=19'b0000000_101110111110;
      15'b001_110110110101 : VALUE=19'b0000000_101110111110;
      15'b001_110110110110 : VALUE=19'b0000000_101110111110;
      15'b001_110110110111 : VALUE=19'b0000000_101110111110;
      15'b001_110110111000 : VALUE=19'b0000000_101110111101;
      15'b001_110110111001 : VALUE=19'b0000000_101110111101;
      15'b001_110110111010 : VALUE=19'b0000000_101110111101;
      15'b001_110110111011 : VALUE=19'b0000000_101110111101;
      15'b001_110110111100 : VALUE=19'b0000000_101110111101;
      15'b001_110110111101 : VALUE=19'b0000000_101110111100;
      15'b001_110110111110 : VALUE=19'b0000000_101110111100;
      15'b001_110110111111 : VALUE=19'b0000000_101110111100;
      15'b001_110111000000 : VALUE=19'b0000000_101110111100;
      15'b001_110111000001 : VALUE=19'b0000000_101110111100;
      15'b001_110111000010 : VALUE=19'b0000000_101110111011;
      15'b001_110111000011 : VALUE=19'b0000000_101110111011;
      15'b001_110111000100 : VALUE=19'b0000000_101110111011;
      15'b001_110111000101 : VALUE=19'b0000000_101110111011;
      15'b001_110111000110 : VALUE=19'b0000000_101110111011;
      15'b001_110111000111 : VALUE=19'b0000000_101110111010;
      15'b001_110111001000 : VALUE=19'b0000000_101110111010;
      15'b001_110111001001 : VALUE=19'b0000000_101110111010;
      15'b001_110111001010 : VALUE=19'b0000000_101110111010;
      15'b001_110111001011 : VALUE=19'b0000000_101110111010;
      15'b001_110111001100 : VALUE=19'b0000000_101110111001;
      15'b001_110111001101 : VALUE=19'b0000000_101110111001;
      15'b001_110111001110 : VALUE=19'b0000000_101110111001;
      15'b001_110111001111 : VALUE=19'b0000000_101110111001;
      15'b001_110111010000 : VALUE=19'b0000000_101110111001;
      15'b001_110111010001 : VALUE=19'b0000000_101110111000;
      15'b001_110111010010 : VALUE=19'b0000000_101110111000;
      15'b001_110111010011 : VALUE=19'b0000000_101110111000;
      15'b001_110111010100 : VALUE=19'b0000000_101110111000;
      15'b001_110111010101 : VALUE=19'b0000000_101110111000;
      15'b001_110111010110 : VALUE=19'b0000000_101110111000;
      15'b001_110111010111 : VALUE=19'b0000000_101110110111;
      15'b001_110111011000 : VALUE=19'b0000000_101110110111;
      15'b001_110111011001 : VALUE=19'b0000000_101110110111;
      15'b001_110111011010 : VALUE=19'b0000000_101110110111;
      15'b001_110111011011 : VALUE=19'b0000000_101110110111;
      15'b001_110111011100 : VALUE=19'b0000000_101110110110;
      15'b001_110111011101 : VALUE=19'b0000000_101110110110;
      15'b001_110111011110 : VALUE=19'b0000000_101110110110;
      15'b001_110111011111 : VALUE=19'b0000000_101110110110;
      15'b001_110111100000 : VALUE=19'b0000000_101110110110;
      15'b001_110111100001 : VALUE=19'b0000000_101110110101;
      15'b001_110111100010 : VALUE=19'b0000000_101110110101;
      15'b001_110111100011 : VALUE=19'b0000000_101110110101;
      15'b001_110111100100 : VALUE=19'b0000000_101110110101;
      15'b001_110111100101 : VALUE=19'b0000000_101110110101;
      15'b001_110111100110 : VALUE=19'b0000000_101110110100;
      15'b001_110111100111 : VALUE=19'b0000000_101110110100;
      15'b001_110111101000 : VALUE=19'b0000000_101110110100;
      15'b001_110111101001 : VALUE=19'b0000000_101110110100;
      15'b001_110111101010 : VALUE=19'b0000000_101110110100;
      15'b001_110111101011 : VALUE=19'b0000000_101110110011;
      15'b001_110111101100 : VALUE=19'b0000000_101110110011;
      15'b001_110111101101 : VALUE=19'b0000000_101110110011;
      15'b001_110111101110 : VALUE=19'b0000000_101110110011;
      15'b001_110111101111 : VALUE=19'b0000000_101110110011;
      15'b001_110111110000 : VALUE=19'b0000000_101110110010;
      15'b001_110111110001 : VALUE=19'b0000000_101110110010;
      15'b001_110111110010 : VALUE=19'b0000000_101110110010;
      15'b001_110111110011 : VALUE=19'b0000000_101110110010;
      15'b001_110111110100 : VALUE=19'b0000000_101110110010;
      15'b001_110111110101 : VALUE=19'b0000000_101110110001;
      15'b001_110111110110 : VALUE=19'b0000000_101110110001;
      15'b001_110111110111 : VALUE=19'b0000000_101110110001;
      15'b001_110111111000 : VALUE=19'b0000000_101110110001;
      15'b001_110111111001 : VALUE=19'b0000000_101110110001;
      15'b001_110111111010 : VALUE=19'b0000000_101110110000;
      15'b001_110111111011 : VALUE=19'b0000000_101110110000;
      15'b001_110111111100 : VALUE=19'b0000000_101110110000;
      15'b001_110111111101 : VALUE=19'b0000000_101110110000;
      15'b001_110111111110 : VALUE=19'b0000000_101110110000;
      15'b001_110111111111 : VALUE=19'b0000000_101110101111;
      15'b001_111000000000 : VALUE=19'b0000000_101110101111;
      15'b001_111000000001 : VALUE=19'b0000000_101110101111;
      15'b001_111000000010 : VALUE=19'b0000000_101110101111;
      15'b001_111000000011 : VALUE=19'b0000000_101110101111;
      15'b001_111000000100 : VALUE=19'b0000000_101110101111;
      15'b001_111000000101 : VALUE=19'b0000000_101110101110;
      15'b001_111000000110 : VALUE=19'b0000000_101110101110;
      15'b001_111000000111 : VALUE=19'b0000000_101110101110;
      15'b001_111000001000 : VALUE=19'b0000000_101110101110;
      15'b001_111000001001 : VALUE=19'b0000000_101110101110;
      15'b001_111000001010 : VALUE=19'b0000000_101110101101;
      15'b001_111000001011 : VALUE=19'b0000000_101110101101;
      15'b001_111000001100 : VALUE=19'b0000000_101110101101;
      15'b001_111000001101 : VALUE=19'b0000000_101110101101;
      15'b001_111000001110 : VALUE=19'b0000000_101110101101;
      15'b001_111000001111 : VALUE=19'b0000000_101110101100;
      15'b001_111000010000 : VALUE=19'b0000000_101110101100;
      15'b001_111000010001 : VALUE=19'b0000000_101110101100;
      15'b001_111000010010 : VALUE=19'b0000000_101110101100;
      15'b001_111000010011 : VALUE=19'b0000000_101110101100;
      15'b001_111000010100 : VALUE=19'b0000000_101110101011;
      15'b001_111000010101 : VALUE=19'b0000000_101110101011;
      15'b001_111000010110 : VALUE=19'b0000000_101110101011;
      15'b001_111000010111 : VALUE=19'b0000000_101110101011;
      15'b001_111000011000 : VALUE=19'b0000000_101110101011;
      15'b001_111000011001 : VALUE=19'b0000000_101110101010;
      15'b001_111000011010 : VALUE=19'b0000000_101110101010;
      15'b001_111000011011 : VALUE=19'b0000000_101110101010;
      15'b001_111000011100 : VALUE=19'b0000000_101110101010;
      15'b001_111000011101 : VALUE=19'b0000000_101110101010;
      15'b001_111000011110 : VALUE=19'b0000000_101110101001;
      15'b001_111000011111 : VALUE=19'b0000000_101110101001;
      15'b001_111000100000 : VALUE=19'b0000000_101110101001;
      15'b001_111000100001 : VALUE=19'b0000000_101110101001;
      15'b001_111000100010 : VALUE=19'b0000000_101110101001;
      15'b001_111000100011 : VALUE=19'b0000000_101110101001;
      15'b001_111000100100 : VALUE=19'b0000000_101110101000;
      15'b001_111000100101 : VALUE=19'b0000000_101110101000;
      15'b001_111000100110 : VALUE=19'b0000000_101110101000;
      15'b001_111000100111 : VALUE=19'b0000000_101110101000;
      15'b001_111000101000 : VALUE=19'b0000000_101110101000;
      15'b001_111000101001 : VALUE=19'b0000000_101110100111;
      15'b001_111000101010 : VALUE=19'b0000000_101110100111;
      15'b001_111000101011 : VALUE=19'b0000000_101110100111;
      15'b001_111000101100 : VALUE=19'b0000000_101110100111;
      15'b001_111000101101 : VALUE=19'b0000000_101110100111;
      15'b001_111000101110 : VALUE=19'b0000000_101110100110;
      15'b001_111000101111 : VALUE=19'b0000000_101110100110;
      15'b001_111000110000 : VALUE=19'b0000000_101110100110;
      15'b001_111000110001 : VALUE=19'b0000000_101110100110;
      15'b001_111000110010 : VALUE=19'b0000000_101110100110;
      15'b001_111000110011 : VALUE=19'b0000000_101110100101;
      15'b001_111000110100 : VALUE=19'b0000000_101110100101;
      15'b001_111000110101 : VALUE=19'b0000000_101110100101;
      15'b001_111000110110 : VALUE=19'b0000000_101110100101;
      15'b001_111000110111 : VALUE=19'b0000000_101110100101;
      15'b001_111000111000 : VALUE=19'b0000000_101110100100;
      15'b001_111000111001 : VALUE=19'b0000000_101110100100;
      15'b001_111000111010 : VALUE=19'b0000000_101110100100;
      15'b001_111000111011 : VALUE=19'b0000000_101110100100;
      15'b001_111000111100 : VALUE=19'b0000000_101110100100;
      15'b001_111000111101 : VALUE=19'b0000000_101110100011;
      15'b001_111000111110 : VALUE=19'b0000000_101110100011;
      15'b001_111000111111 : VALUE=19'b0000000_101110100011;
      15'b001_111001000000 : VALUE=19'b0000000_101110100011;
      15'b001_111001000001 : VALUE=19'b0000000_101110100011;
      15'b001_111001000010 : VALUE=19'b0000000_101110100011;
      15'b001_111001000011 : VALUE=19'b0000000_101110100010;
      15'b001_111001000100 : VALUE=19'b0000000_101110100010;
      15'b001_111001000101 : VALUE=19'b0000000_101110100010;
      15'b001_111001000110 : VALUE=19'b0000000_101110100010;
      15'b001_111001000111 : VALUE=19'b0000000_101110100010;
      15'b001_111001001000 : VALUE=19'b0000000_101110100001;
      15'b001_111001001001 : VALUE=19'b0000000_101110100001;
      15'b001_111001001010 : VALUE=19'b0000000_101110100001;
      15'b001_111001001011 : VALUE=19'b0000000_101110100001;
      15'b001_111001001100 : VALUE=19'b0000000_101110100001;
      15'b001_111001001101 : VALUE=19'b0000000_101110100000;
      15'b001_111001001110 : VALUE=19'b0000000_101110100000;
      15'b001_111001001111 : VALUE=19'b0000000_101110100000;
      15'b001_111001010000 : VALUE=19'b0000000_101110100000;
      15'b001_111001010001 : VALUE=19'b0000000_101110100000;
      15'b001_111001010010 : VALUE=19'b0000000_101110011111;
      15'b001_111001010011 : VALUE=19'b0000000_101110011111;
      15'b001_111001010100 : VALUE=19'b0000000_101110011111;
      15'b001_111001010101 : VALUE=19'b0000000_101110011111;
      15'b001_111001010110 : VALUE=19'b0000000_101110011111;
      15'b001_111001010111 : VALUE=19'b0000000_101110011110;
      15'b001_111001011000 : VALUE=19'b0000000_101110011110;
      15'b001_111001011001 : VALUE=19'b0000000_101110011110;
      15'b001_111001011010 : VALUE=19'b0000000_101110011110;
      15'b001_111001011011 : VALUE=19'b0000000_101110011110;
      15'b001_111001011100 : VALUE=19'b0000000_101110011110;
      15'b001_111001011101 : VALUE=19'b0000000_101110011101;
      15'b001_111001011110 : VALUE=19'b0000000_101110011101;
      15'b001_111001011111 : VALUE=19'b0000000_101110011101;
      15'b001_111001100000 : VALUE=19'b0000000_101110011101;
      15'b001_111001100001 : VALUE=19'b0000000_101110011101;
      15'b001_111001100010 : VALUE=19'b0000000_101110011100;
      15'b001_111001100011 : VALUE=19'b0000000_101110011100;
      15'b001_111001100100 : VALUE=19'b0000000_101110011100;
      15'b001_111001100101 : VALUE=19'b0000000_101110011100;
      15'b001_111001100110 : VALUE=19'b0000000_101110011100;
      15'b001_111001100111 : VALUE=19'b0000000_101110011011;
      15'b001_111001101000 : VALUE=19'b0000000_101110011011;
      15'b001_111001101001 : VALUE=19'b0000000_101110011011;
      15'b001_111001101010 : VALUE=19'b0000000_101110011011;
      15'b001_111001101011 : VALUE=19'b0000000_101110011011;
      15'b001_111001101100 : VALUE=19'b0000000_101110011010;
      15'b001_111001101101 : VALUE=19'b0000000_101110011010;
      15'b001_111001101110 : VALUE=19'b0000000_101110011010;
      15'b001_111001101111 : VALUE=19'b0000000_101110011010;
      15'b001_111001110000 : VALUE=19'b0000000_101110011010;
      15'b001_111001110001 : VALUE=19'b0000000_101110011010;
      15'b001_111001110010 : VALUE=19'b0000000_101110011001;
      15'b001_111001110011 : VALUE=19'b0000000_101110011001;
      15'b001_111001110100 : VALUE=19'b0000000_101110011001;
      15'b001_111001110101 : VALUE=19'b0000000_101110011001;
      15'b001_111001110110 : VALUE=19'b0000000_101110011001;
      15'b001_111001110111 : VALUE=19'b0000000_101110011000;
      15'b001_111001111000 : VALUE=19'b0000000_101110011000;
      15'b001_111001111001 : VALUE=19'b0000000_101110011000;
      15'b001_111001111010 : VALUE=19'b0000000_101110011000;
      15'b001_111001111011 : VALUE=19'b0000000_101110011000;
      15'b001_111001111100 : VALUE=19'b0000000_101110010111;
      15'b001_111001111101 : VALUE=19'b0000000_101110010111;
      15'b001_111001111110 : VALUE=19'b0000000_101110010111;
      15'b001_111001111111 : VALUE=19'b0000000_101110010111;
      15'b001_111010000000 : VALUE=19'b0000000_101110010111;
      15'b001_111010000001 : VALUE=19'b0000000_101110010110;
      15'b001_111010000010 : VALUE=19'b0000000_101110010110;
      15'b001_111010000011 : VALUE=19'b0000000_101110010110;
      15'b001_111010000100 : VALUE=19'b0000000_101110010110;
      15'b001_111010000101 : VALUE=19'b0000000_101110010110;
      15'b001_111010000110 : VALUE=19'b0000000_101110010110;
      15'b001_111010000111 : VALUE=19'b0000000_101110010101;
      15'b001_111010001000 : VALUE=19'b0000000_101110010101;
      15'b001_111010001001 : VALUE=19'b0000000_101110010101;
      15'b001_111010001010 : VALUE=19'b0000000_101110010101;
      15'b001_111010001011 : VALUE=19'b0000000_101110010101;
      15'b001_111010001100 : VALUE=19'b0000000_101110010100;
      15'b001_111010001101 : VALUE=19'b0000000_101110010100;
      15'b001_111010001110 : VALUE=19'b0000000_101110010100;
      15'b001_111010001111 : VALUE=19'b0000000_101110010100;
      15'b001_111010010000 : VALUE=19'b0000000_101110010100;
      15'b001_111010010001 : VALUE=19'b0000000_101110010011;
      15'b001_111010010010 : VALUE=19'b0000000_101110010011;
      15'b001_111010010011 : VALUE=19'b0000000_101110010011;
      15'b001_111010010100 : VALUE=19'b0000000_101110010011;
      15'b001_111010010101 : VALUE=19'b0000000_101110010011;
      15'b001_111010010110 : VALUE=19'b0000000_101110010011;
      15'b001_111010010111 : VALUE=19'b0000000_101110010010;
      15'b001_111010011000 : VALUE=19'b0000000_101110010010;
      15'b001_111010011001 : VALUE=19'b0000000_101110010010;
      15'b001_111010011010 : VALUE=19'b0000000_101110010010;
      15'b001_111010011011 : VALUE=19'b0000000_101110010010;
      15'b001_111010011100 : VALUE=19'b0000000_101110010001;
      15'b001_111010011101 : VALUE=19'b0000000_101110010001;
      15'b001_111010011110 : VALUE=19'b0000000_101110010001;
      15'b001_111010011111 : VALUE=19'b0000000_101110010001;
      15'b001_111010100000 : VALUE=19'b0000000_101110010001;
      15'b001_111010100001 : VALUE=19'b0000000_101110010000;
      15'b001_111010100010 : VALUE=19'b0000000_101110010000;
      15'b001_111010100011 : VALUE=19'b0000000_101110010000;
      15'b001_111010100100 : VALUE=19'b0000000_101110010000;
      15'b001_111010100101 : VALUE=19'b0000000_101110010000;
      15'b001_111010100110 : VALUE=19'b0000000_101110001111;
      15'b001_111010100111 : VALUE=19'b0000000_101110001111;
      15'b001_111010101000 : VALUE=19'b0000000_101110001111;
      15'b001_111010101001 : VALUE=19'b0000000_101110001111;
      15'b001_111010101010 : VALUE=19'b0000000_101110001111;
      15'b001_111010101011 : VALUE=19'b0000000_101110001111;
      15'b001_111010101100 : VALUE=19'b0000000_101110001110;
      15'b001_111010101101 : VALUE=19'b0000000_101110001110;
      15'b001_111010101110 : VALUE=19'b0000000_101110001110;
      15'b001_111010101111 : VALUE=19'b0000000_101110001110;
      15'b001_111010110000 : VALUE=19'b0000000_101110001110;
      15'b001_111010110001 : VALUE=19'b0000000_101110001101;
      15'b001_111010110010 : VALUE=19'b0000000_101110001101;
      15'b001_111010110011 : VALUE=19'b0000000_101110001101;
      15'b001_111010110100 : VALUE=19'b0000000_101110001101;
      15'b001_111010110101 : VALUE=19'b0000000_101110001101;
      15'b001_111010110110 : VALUE=19'b0000000_101110001100;
      15'b001_111010110111 : VALUE=19'b0000000_101110001100;
      15'b001_111010111000 : VALUE=19'b0000000_101110001100;
      15'b001_111010111001 : VALUE=19'b0000000_101110001100;
      15'b001_111010111010 : VALUE=19'b0000000_101110001100;
      15'b001_111010111011 : VALUE=19'b0000000_101110001100;
      15'b001_111010111100 : VALUE=19'b0000000_101110001011;
      15'b001_111010111101 : VALUE=19'b0000000_101110001011;
      15'b001_111010111110 : VALUE=19'b0000000_101110001011;
      15'b001_111010111111 : VALUE=19'b0000000_101110001011;
      15'b001_111011000000 : VALUE=19'b0000000_101110001011;
      15'b001_111011000001 : VALUE=19'b0000000_101110001010;
      15'b001_111011000010 : VALUE=19'b0000000_101110001010;
      15'b001_111011000011 : VALUE=19'b0000000_101110001010;
      15'b001_111011000100 : VALUE=19'b0000000_101110001010;
      15'b001_111011000101 : VALUE=19'b0000000_101110001010;
      15'b001_111011000110 : VALUE=19'b0000000_101110001001;
      15'b001_111011000111 : VALUE=19'b0000000_101110001001;
      15'b001_111011001000 : VALUE=19'b0000000_101110001001;
      15'b001_111011001001 : VALUE=19'b0000000_101110001001;
      15'b001_111011001010 : VALUE=19'b0000000_101110001001;
      15'b001_111011001011 : VALUE=19'b0000000_101110001001;
      15'b001_111011001100 : VALUE=19'b0000000_101110001000;
      15'b001_111011001101 : VALUE=19'b0000000_101110001000;
      15'b001_111011001110 : VALUE=19'b0000000_101110001000;
      15'b001_111011001111 : VALUE=19'b0000000_101110001000;
      15'b001_111011010000 : VALUE=19'b0000000_101110001000;
      15'b001_111011010001 : VALUE=19'b0000000_101110000111;
      15'b001_111011010010 : VALUE=19'b0000000_101110000111;
      15'b001_111011010011 : VALUE=19'b0000000_101110000111;
      15'b001_111011010100 : VALUE=19'b0000000_101110000111;
      15'b001_111011010101 : VALUE=19'b0000000_101110000111;
      15'b001_111011010110 : VALUE=19'b0000000_101110000110;
      15'b001_111011010111 : VALUE=19'b0000000_101110000110;
      15'b001_111011011000 : VALUE=19'b0000000_101110000110;
      15'b001_111011011001 : VALUE=19'b0000000_101110000110;
      15'b001_111011011010 : VALUE=19'b0000000_101110000110;
      15'b001_111011011011 : VALUE=19'b0000000_101110000110;
      15'b001_111011011100 : VALUE=19'b0000000_101110000101;
      15'b001_111011011101 : VALUE=19'b0000000_101110000101;
      15'b001_111011011110 : VALUE=19'b0000000_101110000101;
      15'b001_111011011111 : VALUE=19'b0000000_101110000101;
      15'b001_111011100000 : VALUE=19'b0000000_101110000101;
      15'b001_111011100001 : VALUE=19'b0000000_101110000100;
      15'b001_111011100010 : VALUE=19'b0000000_101110000100;
      15'b001_111011100011 : VALUE=19'b0000000_101110000100;
      15'b001_111011100100 : VALUE=19'b0000000_101110000100;
      15'b001_111011100101 : VALUE=19'b0000000_101110000100;
      15'b001_111011100110 : VALUE=19'b0000000_101110000011;
      15'b001_111011100111 : VALUE=19'b0000000_101110000011;
      15'b001_111011101000 : VALUE=19'b0000000_101110000011;
      15'b001_111011101001 : VALUE=19'b0000000_101110000011;
      15'b001_111011101010 : VALUE=19'b0000000_101110000011;
      15'b001_111011101011 : VALUE=19'b0000000_101110000011;
      15'b001_111011101100 : VALUE=19'b0000000_101110000010;
      15'b001_111011101101 : VALUE=19'b0000000_101110000010;
      15'b001_111011101110 : VALUE=19'b0000000_101110000010;
      15'b001_111011101111 : VALUE=19'b0000000_101110000010;
      15'b001_111011110000 : VALUE=19'b0000000_101110000010;
      15'b001_111011110001 : VALUE=19'b0000000_101110000001;
      15'b001_111011110010 : VALUE=19'b0000000_101110000001;
      15'b001_111011110011 : VALUE=19'b0000000_101110000001;
      15'b001_111011110100 : VALUE=19'b0000000_101110000001;
      15'b001_111011110101 : VALUE=19'b0000000_101110000001;
      15'b001_111011110110 : VALUE=19'b0000000_101110000001;
      15'b001_111011110111 : VALUE=19'b0000000_101110000000;
      15'b001_111011111000 : VALUE=19'b0000000_101110000000;
      15'b001_111011111001 : VALUE=19'b0000000_101110000000;
      15'b001_111011111010 : VALUE=19'b0000000_101110000000;
      15'b001_111011111011 : VALUE=19'b0000000_101110000000;
      15'b001_111011111100 : VALUE=19'b0000000_101101111111;
      15'b001_111011111101 : VALUE=19'b0000000_101101111111;
      15'b001_111011111110 : VALUE=19'b0000000_101101111111;
      15'b001_111011111111 : VALUE=19'b0000000_101101111111;
      15'b001_111100000000 : VALUE=19'b0000000_101101111111;
      15'b001_111100000001 : VALUE=19'b0000000_101101111110;
      15'b001_111100000010 : VALUE=19'b0000000_101101111110;
      15'b001_111100000011 : VALUE=19'b0000000_101101111110;
      15'b001_111100000100 : VALUE=19'b0000000_101101111110;
      15'b001_111100000101 : VALUE=19'b0000000_101101111110;
      15'b001_111100000110 : VALUE=19'b0000000_101101111110;
      15'b001_111100000111 : VALUE=19'b0000000_101101111101;
      15'b001_111100001000 : VALUE=19'b0000000_101101111101;
      15'b001_111100001001 : VALUE=19'b0000000_101101111101;
      15'b001_111100001010 : VALUE=19'b0000000_101101111101;
      15'b001_111100001011 : VALUE=19'b0000000_101101111101;
      15'b001_111100001100 : VALUE=19'b0000000_101101111100;
      15'b001_111100001101 : VALUE=19'b0000000_101101111100;
      15'b001_111100001110 : VALUE=19'b0000000_101101111100;
      15'b001_111100001111 : VALUE=19'b0000000_101101111100;
      15'b001_111100010000 : VALUE=19'b0000000_101101111100;
      15'b001_111100010001 : VALUE=19'b0000000_101101111100;
      15'b001_111100010010 : VALUE=19'b0000000_101101111011;
      15'b001_111100010011 : VALUE=19'b0000000_101101111011;
      15'b001_111100010100 : VALUE=19'b0000000_101101111011;
      15'b001_111100010101 : VALUE=19'b0000000_101101111011;
      15'b001_111100010110 : VALUE=19'b0000000_101101111011;
      15'b001_111100010111 : VALUE=19'b0000000_101101111010;
      15'b001_111100011000 : VALUE=19'b0000000_101101111010;
      15'b001_111100011001 : VALUE=19'b0000000_101101111010;
      15'b001_111100011010 : VALUE=19'b0000000_101101111010;
      15'b001_111100011011 : VALUE=19'b0000000_101101111010;
      15'b001_111100011100 : VALUE=19'b0000000_101101111001;
      15'b001_111100011101 : VALUE=19'b0000000_101101111001;
      15'b001_111100011110 : VALUE=19'b0000000_101101111001;
      15'b001_111100011111 : VALUE=19'b0000000_101101111001;
      15'b001_111100100000 : VALUE=19'b0000000_101101111001;
      15'b001_111100100001 : VALUE=19'b0000000_101101111001;
      15'b001_111100100010 : VALUE=19'b0000000_101101111000;
      15'b001_111100100011 : VALUE=19'b0000000_101101111000;
      15'b001_111100100100 : VALUE=19'b0000000_101101111000;
      15'b001_111100100101 : VALUE=19'b0000000_101101111000;
      15'b001_111100100110 : VALUE=19'b0000000_101101111000;
      15'b001_111100100111 : VALUE=19'b0000000_101101110111;
      15'b001_111100101000 : VALUE=19'b0000000_101101110111;
      15'b001_111100101001 : VALUE=19'b0000000_101101110111;
      15'b001_111100101010 : VALUE=19'b0000000_101101110111;
      15'b001_111100101011 : VALUE=19'b0000000_101101110111;
      15'b001_111100101100 : VALUE=19'b0000000_101101110111;
      15'b001_111100101101 : VALUE=19'b0000000_101101110110;
      15'b001_111100101110 : VALUE=19'b0000000_101101110110;
      15'b001_111100101111 : VALUE=19'b0000000_101101110110;
      15'b001_111100110000 : VALUE=19'b0000000_101101110110;
      15'b001_111100110001 : VALUE=19'b0000000_101101110110;
      15'b001_111100110010 : VALUE=19'b0000000_101101110101;
      15'b001_111100110011 : VALUE=19'b0000000_101101110101;
      15'b001_111100110100 : VALUE=19'b0000000_101101110101;
      15'b001_111100110101 : VALUE=19'b0000000_101101110101;
      15'b001_111100110110 : VALUE=19'b0000000_101101110101;
      15'b001_111100110111 : VALUE=19'b0000000_101101110101;
      15'b001_111100111000 : VALUE=19'b0000000_101101110100;
      15'b001_111100111001 : VALUE=19'b0000000_101101110100;
      15'b001_111100111010 : VALUE=19'b0000000_101101110100;
      15'b001_111100111011 : VALUE=19'b0000000_101101110100;
      15'b001_111100111100 : VALUE=19'b0000000_101101110100;
      15'b001_111100111101 : VALUE=19'b0000000_101101110011;
      15'b001_111100111110 : VALUE=19'b0000000_101101110011;
      15'b001_111100111111 : VALUE=19'b0000000_101101110011;
      15'b001_111101000000 : VALUE=19'b0000000_101101110011;
      15'b001_111101000001 : VALUE=19'b0000000_101101110011;
      15'b001_111101000010 : VALUE=19'b0000000_101101110010;
      15'b001_111101000011 : VALUE=19'b0000000_101101110010;
      15'b001_111101000100 : VALUE=19'b0000000_101101110010;
      15'b001_111101000101 : VALUE=19'b0000000_101101110010;
      15'b001_111101000110 : VALUE=19'b0000000_101101110010;
      15'b001_111101000111 : VALUE=19'b0000000_101101110010;
      15'b001_111101001000 : VALUE=19'b0000000_101101110001;
      15'b001_111101001001 : VALUE=19'b0000000_101101110001;
      15'b001_111101001010 : VALUE=19'b0000000_101101110001;
      15'b001_111101001011 : VALUE=19'b0000000_101101110001;
      15'b001_111101001100 : VALUE=19'b0000000_101101110001;
      15'b001_111101001101 : VALUE=19'b0000000_101101110000;
      15'b001_111101001110 : VALUE=19'b0000000_101101110000;
      15'b001_111101001111 : VALUE=19'b0000000_101101110000;
      15'b001_111101010000 : VALUE=19'b0000000_101101110000;
      15'b001_111101010001 : VALUE=19'b0000000_101101110000;
      15'b001_111101010010 : VALUE=19'b0000000_101101110000;
      15'b001_111101010011 : VALUE=19'b0000000_101101101111;
      15'b001_111101010100 : VALUE=19'b0000000_101101101111;
      15'b001_111101010101 : VALUE=19'b0000000_101101101111;
      15'b001_111101010110 : VALUE=19'b0000000_101101101111;
      15'b001_111101010111 : VALUE=19'b0000000_101101101111;
      15'b001_111101011000 : VALUE=19'b0000000_101101101110;
      15'b001_111101011001 : VALUE=19'b0000000_101101101110;
      15'b001_111101011010 : VALUE=19'b0000000_101101101110;
      15'b001_111101011011 : VALUE=19'b0000000_101101101110;
      15'b001_111101011100 : VALUE=19'b0000000_101101101110;
      15'b001_111101011101 : VALUE=19'b0000000_101101101110;
      15'b001_111101011110 : VALUE=19'b0000000_101101101101;
      15'b001_111101011111 : VALUE=19'b0000000_101101101101;
      15'b001_111101100000 : VALUE=19'b0000000_101101101101;
      15'b001_111101100001 : VALUE=19'b0000000_101101101101;
      15'b001_111101100010 : VALUE=19'b0000000_101101101101;
      15'b001_111101100011 : VALUE=19'b0000000_101101101100;
      15'b001_111101100100 : VALUE=19'b0000000_101101101100;
      15'b001_111101100101 : VALUE=19'b0000000_101101101100;
      15'b001_111101100110 : VALUE=19'b0000000_101101101100;
      15'b001_111101100111 : VALUE=19'b0000000_101101101100;
      15'b001_111101101000 : VALUE=19'b0000000_101101101100;
      15'b001_111101101001 : VALUE=19'b0000000_101101101011;
      15'b001_111101101010 : VALUE=19'b0000000_101101101011;
      15'b001_111101101011 : VALUE=19'b0000000_101101101011;
      15'b001_111101101100 : VALUE=19'b0000000_101101101011;
      15'b001_111101101101 : VALUE=19'b0000000_101101101011;
      15'b001_111101101110 : VALUE=19'b0000000_101101101010;
      15'b001_111101101111 : VALUE=19'b0000000_101101101010;
      15'b001_111101110000 : VALUE=19'b0000000_101101101010;
      15'b001_111101110001 : VALUE=19'b0000000_101101101010;
      15'b001_111101110010 : VALUE=19'b0000000_101101101010;
      15'b001_111101110011 : VALUE=19'b0000000_101101101010;
      15'b001_111101110100 : VALUE=19'b0000000_101101101001;
      15'b001_111101110101 : VALUE=19'b0000000_101101101001;
      15'b001_111101110110 : VALUE=19'b0000000_101101101001;
      15'b001_111101110111 : VALUE=19'b0000000_101101101001;
      15'b001_111101111000 : VALUE=19'b0000000_101101101001;
      15'b001_111101111001 : VALUE=19'b0000000_101101101000;
      15'b001_111101111010 : VALUE=19'b0000000_101101101000;
      15'b001_111101111011 : VALUE=19'b0000000_101101101000;
      15'b001_111101111100 : VALUE=19'b0000000_101101101000;
      15'b001_111101111101 : VALUE=19'b0000000_101101101000;
      15'b001_111101111110 : VALUE=19'b0000000_101101101000;
      15'b001_111101111111 : VALUE=19'b0000000_101101100111;
      15'b001_111110000000 : VALUE=19'b0000000_101101100111;
      15'b001_111110000001 : VALUE=19'b0000000_101101100111;
      15'b001_111110000010 : VALUE=19'b0000000_101101100111;
      15'b001_111110000011 : VALUE=19'b0000000_101101100111;
      15'b001_111110000100 : VALUE=19'b0000000_101101100110;
      15'b001_111110000101 : VALUE=19'b0000000_101101100110;
      15'b001_111110000110 : VALUE=19'b0000000_101101100110;
      15'b001_111110000111 : VALUE=19'b0000000_101101100110;
      15'b001_111110001000 : VALUE=19'b0000000_101101100110;
      15'b001_111110001001 : VALUE=19'b0000000_101101100110;
      15'b001_111110001010 : VALUE=19'b0000000_101101100101;
      15'b001_111110001011 : VALUE=19'b0000000_101101100101;
      15'b001_111110001100 : VALUE=19'b0000000_101101100101;
      15'b001_111110001101 : VALUE=19'b0000000_101101100101;
      15'b001_111110001110 : VALUE=19'b0000000_101101100101;
      15'b001_111110001111 : VALUE=19'b0000000_101101100100;
      15'b001_111110010000 : VALUE=19'b0000000_101101100100;
      15'b001_111110010001 : VALUE=19'b0000000_101101100100;
      15'b001_111110010010 : VALUE=19'b0000000_101101100100;
      15'b001_111110010011 : VALUE=19'b0000000_101101100100;
      15'b001_111110010100 : VALUE=19'b0000000_101101100100;
      15'b001_111110010101 : VALUE=19'b0000000_101101100011;
      15'b001_111110010110 : VALUE=19'b0000000_101101100011;
      15'b001_111110010111 : VALUE=19'b0000000_101101100011;
      15'b001_111110011000 : VALUE=19'b0000000_101101100011;
      15'b001_111110011001 : VALUE=19'b0000000_101101100011;
      15'b001_111110011010 : VALUE=19'b0000000_101101100011;
      15'b001_111110011011 : VALUE=19'b0000000_101101100010;
      15'b001_111110011100 : VALUE=19'b0000000_101101100010;
      15'b001_111110011101 : VALUE=19'b0000000_101101100010;
      15'b001_111110011110 : VALUE=19'b0000000_101101100010;
      15'b001_111110011111 : VALUE=19'b0000000_101101100010;
      15'b001_111110100000 : VALUE=19'b0000000_101101100001;
      15'b001_111110100001 : VALUE=19'b0000000_101101100001;
      15'b001_111110100010 : VALUE=19'b0000000_101101100001;
      15'b001_111110100011 : VALUE=19'b0000000_101101100001;
      15'b001_111110100100 : VALUE=19'b0000000_101101100001;
      15'b001_111110100101 : VALUE=19'b0000000_101101100001;
      15'b001_111110100110 : VALUE=19'b0000000_101101100000;
      15'b001_111110100111 : VALUE=19'b0000000_101101100000;
      15'b001_111110101000 : VALUE=19'b0000000_101101100000;
      15'b001_111110101001 : VALUE=19'b0000000_101101100000;
      15'b001_111110101010 : VALUE=19'b0000000_101101100000;
      15'b001_111110101011 : VALUE=19'b0000000_101101011111;
      15'b001_111110101100 : VALUE=19'b0000000_101101011111;
      15'b001_111110101101 : VALUE=19'b0000000_101101011111;
      15'b001_111110101110 : VALUE=19'b0000000_101101011111;
      15'b001_111110101111 : VALUE=19'b0000000_101101011111;
      15'b001_111110110000 : VALUE=19'b0000000_101101011111;
      15'b001_111110110001 : VALUE=19'b0000000_101101011110;
      15'b001_111110110010 : VALUE=19'b0000000_101101011110;
      15'b001_111110110011 : VALUE=19'b0000000_101101011110;
      15'b001_111110110100 : VALUE=19'b0000000_101101011110;
      15'b001_111110110101 : VALUE=19'b0000000_101101011110;
      15'b001_111110110110 : VALUE=19'b0000000_101101011101;
      15'b001_111110110111 : VALUE=19'b0000000_101101011101;
      15'b001_111110111000 : VALUE=19'b0000000_101101011101;
      15'b001_111110111001 : VALUE=19'b0000000_101101011101;
      15'b001_111110111010 : VALUE=19'b0000000_101101011101;
      15'b001_111110111011 : VALUE=19'b0000000_101101011101;
      15'b001_111110111100 : VALUE=19'b0000000_101101011100;
      15'b001_111110111101 : VALUE=19'b0000000_101101011100;
      15'b001_111110111110 : VALUE=19'b0000000_101101011100;
      15'b001_111110111111 : VALUE=19'b0000000_101101011100;
      15'b001_111111000000 : VALUE=19'b0000000_101101011100;
      15'b001_111111000001 : VALUE=19'b0000000_101101011100;
      15'b001_111111000010 : VALUE=19'b0000000_101101011011;
      15'b001_111111000011 : VALUE=19'b0000000_101101011011;
      15'b001_111111000100 : VALUE=19'b0000000_101101011011;
      15'b001_111111000101 : VALUE=19'b0000000_101101011011;
      15'b001_111111000110 : VALUE=19'b0000000_101101011011;
      15'b001_111111000111 : VALUE=19'b0000000_101101011010;
      15'b001_111111001000 : VALUE=19'b0000000_101101011010;
      15'b001_111111001001 : VALUE=19'b0000000_101101011010;
      15'b001_111111001010 : VALUE=19'b0000000_101101011010;
      15'b001_111111001011 : VALUE=19'b0000000_101101011010;
      15'b001_111111001100 : VALUE=19'b0000000_101101011010;
      15'b001_111111001101 : VALUE=19'b0000000_101101011001;
      15'b001_111111001110 : VALUE=19'b0000000_101101011001;
      15'b001_111111001111 : VALUE=19'b0000000_101101011001;
      15'b001_111111010000 : VALUE=19'b0000000_101101011001;
      15'b001_111111010001 : VALUE=19'b0000000_101101011001;
      15'b001_111111010010 : VALUE=19'b0000000_101101011000;
      15'b001_111111010011 : VALUE=19'b0000000_101101011000;
      15'b001_111111010100 : VALUE=19'b0000000_101101011000;
      15'b001_111111010101 : VALUE=19'b0000000_101101011000;
      15'b001_111111010110 : VALUE=19'b0000000_101101011000;
      15'b001_111111010111 : VALUE=19'b0000000_101101011000;
      15'b001_111111011000 : VALUE=19'b0000000_101101010111;
      15'b001_111111011001 : VALUE=19'b0000000_101101010111;
      15'b001_111111011010 : VALUE=19'b0000000_101101010111;
      15'b001_111111011011 : VALUE=19'b0000000_101101010111;
      15'b001_111111011100 : VALUE=19'b0000000_101101010111;
      15'b001_111111011101 : VALUE=19'b0000000_101101010111;
      15'b001_111111011110 : VALUE=19'b0000000_101101010110;
      15'b001_111111011111 : VALUE=19'b0000000_101101010110;
      15'b001_111111100000 : VALUE=19'b0000000_101101010110;
      15'b001_111111100001 : VALUE=19'b0000000_101101010110;
      15'b001_111111100010 : VALUE=19'b0000000_101101010110;
      15'b001_111111100011 : VALUE=19'b0000000_101101010101;
      15'b001_111111100100 : VALUE=19'b0000000_101101010101;
      15'b001_111111100101 : VALUE=19'b0000000_101101010101;
      15'b001_111111100110 : VALUE=19'b0000000_101101010101;
      15'b001_111111100111 : VALUE=19'b0000000_101101010101;
      15'b001_111111101000 : VALUE=19'b0000000_101101010101;
      15'b001_111111101001 : VALUE=19'b0000000_101101010100;
      15'b001_111111101010 : VALUE=19'b0000000_101101010100;
      15'b001_111111101011 : VALUE=19'b0000000_101101010100;
      15'b001_111111101100 : VALUE=19'b0000000_101101010100;
      15'b001_111111101101 : VALUE=19'b0000000_101101010100;
      15'b001_111111101110 : VALUE=19'b0000000_101101010011;
      15'b001_111111101111 : VALUE=19'b0000000_101101010011;
      15'b001_111111110000 : VALUE=19'b0000000_101101010011;
      15'b001_111111110001 : VALUE=19'b0000000_101101010011;
      15'b001_111111110010 : VALUE=19'b0000000_101101010011;
      15'b001_111111110011 : VALUE=19'b0000000_101101010011;
      15'b001_111111110100 : VALUE=19'b0000000_101101010010;
      15'b001_111111110101 : VALUE=19'b0000000_101101010010;
      15'b001_111111110110 : VALUE=19'b0000000_101101010010;
      15'b001_111111110111 : VALUE=19'b0000000_101101010010;
      15'b001_111111111000 : VALUE=19'b0000000_101101010010;
      15'b001_111111111001 : VALUE=19'b0000000_101101010010;
      15'b001_111111111010 : VALUE=19'b0000000_101101010001;
      15'b001_111111111011 : VALUE=19'b0000000_101101010001;
      15'b001_111111111100 : VALUE=19'b0000000_101101010001;
      15'b001_111111111101 : VALUE=19'b0000000_101101010001;
      15'b001_111111111110 : VALUE=19'b0000000_101101010001;
      15'b001_111111111111 : VALUE=19'b0000000_101101010000;
      15'b010_000000000000 : VALUE=19'b0000000_101101010000;
      15'b010_000000000001 : VALUE=19'b0000000_101101010000;
      15'b010_000000000010 : VALUE=19'b0000000_101101010000;
      15'b010_000000000011 : VALUE=19'b0000000_101101010000;
      15'b010_000000000100 : VALUE=19'b0000000_101101010000;
      15'b010_000000000101 : VALUE=19'b0000000_101101001111;
      15'b010_000000000110 : VALUE=19'b0000000_101101001111;
      15'b010_000000000111 : VALUE=19'b0000000_101101001111;
      15'b010_000000001000 : VALUE=19'b0000000_101101001111;
      15'b010_000000001001 : VALUE=19'b0000000_101101001111;
      15'b010_000000001010 : VALUE=19'b0000000_101101001111;
      15'b010_000000001011 : VALUE=19'b0000000_101101001110;
      15'b010_000000001100 : VALUE=19'b0000000_101101001110;
      15'b010_000000001101 : VALUE=19'b0000000_101101001110;
      15'b010_000000001110 : VALUE=19'b0000000_101101001110;
      15'b010_000000001111 : VALUE=19'b0000000_101101001110;
      15'b010_000000010000 : VALUE=19'b0000000_101101001101;
      15'b010_000000010001 : VALUE=19'b0000000_101101001101;
      15'b010_000000010010 : VALUE=19'b0000000_101101001101;
      15'b010_000000010011 : VALUE=19'b0000000_101101001101;
      15'b010_000000010100 : VALUE=19'b0000000_101101001101;
      15'b010_000000010101 : VALUE=19'b0000000_101101001101;
      15'b010_000000010110 : VALUE=19'b0000000_101101001100;
      15'b010_000000010111 : VALUE=19'b0000000_101101001100;
      15'b010_000000011000 : VALUE=19'b0000000_101101001100;
      15'b010_000000011001 : VALUE=19'b0000000_101101001100;
      15'b010_000000011010 : VALUE=19'b0000000_101101001100;
      15'b010_000000011011 : VALUE=19'b0000000_101101001100;
      15'b010_000000011100 : VALUE=19'b0000000_101101001011;
      15'b010_000000011101 : VALUE=19'b0000000_101101001011;
      15'b010_000000011110 : VALUE=19'b0000000_101101001011;
      15'b010_000000011111 : VALUE=19'b0000000_101101001011;
      15'b010_000000100000 : VALUE=19'b0000000_101101001011;
      15'b010_000000100001 : VALUE=19'b0000000_101101001010;
      15'b010_000000100010 : VALUE=19'b0000000_101101001010;
      15'b010_000000100011 : VALUE=19'b0000000_101101001010;
      15'b010_000000100100 : VALUE=19'b0000000_101101001010;
      15'b010_000000100101 : VALUE=19'b0000000_101101001010;
      15'b010_000000100110 : VALUE=19'b0000000_101101001010;
      15'b010_000000100111 : VALUE=19'b0000000_101101001001;
      15'b010_000000101000 : VALUE=19'b0000000_101101001001;
      15'b010_000000101001 : VALUE=19'b0000000_101101001001;
      15'b010_000000101010 : VALUE=19'b0000000_101101001001;
      15'b010_000000101011 : VALUE=19'b0000000_101101001001;
      15'b010_000000101100 : VALUE=19'b0000000_101101001001;
      15'b010_000000101101 : VALUE=19'b0000000_101101001000;
      15'b010_000000101110 : VALUE=19'b0000000_101101001000;
      15'b010_000000101111 : VALUE=19'b0000000_101101001000;
      15'b010_000000110000 : VALUE=19'b0000000_101101001000;
      15'b010_000000110001 : VALUE=19'b0000000_101101001000;
      15'b010_000000110010 : VALUE=19'b0000000_101101001000;
      15'b010_000000110011 : VALUE=19'b0000000_101101000111;
      15'b010_000000110100 : VALUE=19'b0000000_101101000111;
      15'b010_000000110101 : VALUE=19'b0000000_101101000111;
      15'b010_000000110110 : VALUE=19'b0000000_101101000111;
      15'b010_000000110111 : VALUE=19'b0000000_101101000111;
      15'b010_000000111000 : VALUE=19'b0000000_101101000110;
      15'b010_000000111001 : VALUE=19'b0000000_101101000110;
      15'b010_000000111010 : VALUE=19'b0000000_101101000110;
      15'b010_000000111011 : VALUE=19'b0000000_101101000110;
      15'b010_000000111100 : VALUE=19'b0000000_101101000110;
      15'b010_000000111101 : VALUE=19'b0000000_101101000110;
      15'b010_000000111110 : VALUE=19'b0000000_101101000101;
      15'b010_000000111111 : VALUE=19'b0000000_101101000101;
      15'b010_000001000000 : VALUE=19'b0000000_101101000101;
      15'b010_000001000001 : VALUE=19'b0000000_101101000101;
      15'b010_000001000010 : VALUE=19'b0000000_101101000101;
      15'b010_000001000011 : VALUE=19'b0000000_101101000101;
      15'b010_000001000100 : VALUE=19'b0000000_101101000100;
      15'b010_000001000101 : VALUE=19'b0000000_101101000100;
      15'b010_000001000110 : VALUE=19'b0000000_101101000100;
      15'b010_000001000111 : VALUE=19'b0000000_101101000100;
      15'b010_000001001000 : VALUE=19'b0000000_101101000100;
      15'b010_000001001001 : VALUE=19'b0000000_101101000011;
      15'b010_000001001010 : VALUE=19'b0000000_101101000011;
      15'b010_000001001011 : VALUE=19'b0000000_101101000011;
      15'b010_000001001100 : VALUE=19'b0000000_101101000011;
      15'b010_000001001101 : VALUE=19'b0000000_101101000011;
      15'b010_000001001110 : VALUE=19'b0000000_101101000011;
      15'b010_000001001111 : VALUE=19'b0000000_101101000010;
      15'b010_000001010000 : VALUE=19'b0000000_101101000010;
      15'b010_000001010001 : VALUE=19'b0000000_101101000010;
      15'b010_000001010010 : VALUE=19'b0000000_101101000010;
      15'b010_000001010011 : VALUE=19'b0000000_101101000010;
      15'b010_000001010100 : VALUE=19'b0000000_101101000010;
      15'b010_000001010101 : VALUE=19'b0000000_101101000001;
      15'b010_000001010110 : VALUE=19'b0000000_101101000001;
      15'b010_000001010111 : VALUE=19'b0000000_101101000001;
      15'b010_000001011000 : VALUE=19'b0000000_101101000001;
      15'b010_000001011001 : VALUE=19'b0000000_101101000001;
      15'b010_000001011010 : VALUE=19'b0000000_101101000001;
      15'b010_000001011011 : VALUE=19'b0000000_101101000000;
      15'b010_000001011100 : VALUE=19'b0000000_101101000000;
      15'b010_000001011101 : VALUE=19'b0000000_101101000000;
      15'b010_000001011110 : VALUE=19'b0000000_101101000000;
      15'b010_000001011111 : VALUE=19'b0000000_101101000000;
      15'b010_000001100000 : VALUE=19'b0000000_101100111111;
      15'b010_000001100001 : VALUE=19'b0000000_101100111111;
      15'b010_000001100010 : VALUE=19'b0000000_101100111111;
      15'b010_000001100011 : VALUE=19'b0000000_101100111111;
      15'b010_000001100100 : VALUE=19'b0000000_101100111111;
      15'b010_000001100101 : VALUE=19'b0000000_101100111111;
      15'b010_000001100110 : VALUE=19'b0000000_101100111110;
      15'b010_000001100111 : VALUE=19'b0000000_101100111110;
      15'b010_000001101000 : VALUE=19'b0000000_101100111110;
      15'b010_000001101001 : VALUE=19'b0000000_101100111110;
      15'b010_000001101010 : VALUE=19'b0000000_101100111110;
      15'b010_000001101011 : VALUE=19'b0000000_101100111110;
      15'b010_000001101100 : VALUE=19'b0000000_101100111101;
      15'b010_000001101101 : VALUE=19'b0000000_101100111101;
      15'b010_000001101110 : VALUE=19'b0000000_101100111101;
      15'b010_000001101111 : VALUE=19'b0000000_101100111101;
      15'b010_000001110000 : VALUE=19'b0000000_101100111101;
      15'b010_000001110001 : VALUE=19'b0000000_101100111101;
      15'b010_000001110010 : VALUE=19'b0000000_101100111100;
      15'b010_000001110011 : VALUE=19'b0000000_101100111100;
      15'b010_000001110100 : VALUE=19'b0000000_101100111100;
      15'b010_000001110101 : VALUE=19'b0000000_101100111100;
      15'b010_000001110110 : VALUE=19'b0000000_101100111100;
      15'b010_000001110111 : VALUE=19'b0000000_101100111011;
      15'b010_000001111000 : VALUE=19'b0000000_101100111011;
      15'b010_000001111001 : VALUE=19'b0000000_101100111011;
      15'b010_000001111010 : VALUE=19'b0000000_101100111011;
      15'b010_000001111011 : VALUE=19'b0000000_101100111011;
      15'b010_000001111100 : VALUE=19'b0000000_101100111011;
      15'b010_000001111101 : VALUE=19'b0000000_101100111010;
      15'b010_000001111110 : VALUE=19'b0000000_101100111010;
      15'b010_000001111111 : VALUE=19'b0000000_101100111010;
      15'b010_000010000000 : VALUE=19'b0000000_101100111010;
      15'b010_000010000001 : VALUE=19'b0000000_101100111010;
      15'b010_000010000010 : VALUE=19'b0000000_101100111010;
      15'b010_000010000011 : VALUE=19'b0000000_101100111001;
      15'b010_000010000100 : VALUE=19'b0000000_101100111001;
      15'b010_000010000101 : VALUE=19'b0000000_101100111001;
      15'b010_000010000110 : VALUE=19'b0000000_101100111001;
      15'b010_000010000111 : VALUE=19'b0000000_101100111001;
      15'b010_000010001000 : VALUE=19'b0000000_101100111001;
      15'b010_000010001001 : VALUE=19'b0000000_101100111000;
      15'b010_000010001010 : VALUE=19'b0000000_101100111000;
      15'b010_000010001011 : VALUE=19'b0000000_101100111000;
      15'b010_000010001100 : VALUE=19'b0000000_101100111000;
      15'b010_000010001101 : VALUE=19'b0000000_101100111000;
      15'b010_000010001110 : VALUE=19'b0000000_101100111000;
      15'b010_000010001111 : VALUE=19'b0000000_101100110111;
      15'b010_000010010000 : VALUE=19'b0000000_101100110111;
      15'b010_000010010001 : VALUE=19'b0000000_101100110111;
      15'b010_000010010010 : VALUE=19'b0000000_101100110111;
      15'b010_000010010011 : VALUE=19'b0000000_101100110111;
      15'b010_000010010100 : VALUE=19'b0000000_101100110110;
      15'b010_000010010101 : VALUE=19'b0000000_101100110110;
      15'b010_000010010110 : VALUE=19'b0000000_101100110110;
      15'b010_000010010111 : VALUE=19'b0000000_101100110110;
      15'b010_000010011000 : VALUE=19'b0000000_101100110110;
      15'b010_000010011001 : VALUE=19'b0000000_101100110110;
      15'b010_000010011010 : VALUE=19'b0000000_101100110101;
      15'b010_000010011011 : VALUE=19'b0000000_101100110101;
      15'b010_000010011100 : VALUE=19'b0000000_101100110101;
      15'b010_000010011101 : VALUE=19'b0000000_101100110101;
      15'b010_000010011110 : VALUE=19'b0000000_101100110101;
      15'b010_000010011111 : VALUE=19'b0000000_101100110101;
      15'b010_000010100000 : VALUE=19'b0000000_101100110100;
      15'b010_000010100001 : VALUE=19'b0000000_101100110100;
      15'b010_000010100010 : VALUE=19'b0000000_101100110100;
      15'b010_000010100011 : VALUE=19'b0000000_101100110100;
      15'b010_000010100100 : VALUE=19'b0000000_101100110100;
      15'b010_000010100101 : VALUE=19'b0000000_101100110100;
      15'b010_000010100110 : VALUE=19'b0000000_101100110011;
      15'b010_000010100111 : VALUE=19'b0000000_101100110011;
      15'b010_000010101000 : VALUE=19'b0000000_101100110011;
      15'b010_000010101001 : VALUE=19'b0000000_101100110011;
      15'b010_000010101010 : VALUE=19'b0000000_101100110011;
      15'b010_000010101011 : VALUE=19'b0000000_101100110011;
      15'b010_000010101100 : VALUE=19'b0000000_101100110010;
      15'b010_000010101101 : VALUE=19'b0000000_101100110010;
      15'b010_000010101110 : VALUE=19'b0000000_101100110010;
      15'b010_000010101111 : VALUE=19'b0000000_101100110010;
      15'b010_000010110000 : VALUE=19'b0000000_101100110010;
      15'b010_000010110001 : VALUE=19'b0000000_101100110010;
      15'b010_000010110010 : VALUE=19'b0000000_101100110001;
      15'b010_000010110011 : VALUE=19'b0000000_101100110001;
      15'b010_000010110100 : VALUE=19'b0000000_101100110001;
      15'b010_000010110101 : VALUE=19'b0000000_101100110001;
      15'b010_000010110110 : VALUE=19'b0000000_101100110001;
      15'b010_000010110111 : VALUE=19'b0000000_101100110000;
      15'b010_000010111000 : VALUE=19'b0000000_101100110000;
      15'b010_000010111001 : VALUE=19'b0000000_101100110000;
      15'b010_000010111010 : VALUE=19'b0000000_101100110000;
      15'b010_000010111011 : VALUE=19'b0000000_101100110000;
      15'b010_000010111100 : VALUE=19'b0000000_101100110000;
      15'b010_000010111101 : VALUE=19'b0000000_101100101111;
      15'b010_000010111110 : VALUE=19'b0000000_101100101111;
      15'b010_000010111111 : VALUE=19'b0000000_101100101111;
      15'b010_000011000000 : VALUE=19'b0000000_101100101111;
      15'b010_000011000001 : VALUE=19'b0000000_101100101111;
      15'b010_000011000010 : VALUE=19'b0000000_101100101111;
      15'b010_000011000011 : VALUE=19'b0000000_101100101110;
      15'b010_000011000100 : VALUE=19'b0000000_101100101110;
      15'b010_000011000101 : VALUE=19'b0000000_101100101110;
      15'b010_000011000110 : VALUE=19'b0000000_101100101110;
      15'b010_000011000111 : VALUE=19'b0000000_101100101110;
      15'b010_000011001000 : VALUE=19'b0000000_101100101110;
      15'b010_000011001001 : VALUE=19'b0000000_101100101101;
      15'b010_000011001010 : VALUE=19'b0000000_101100101101;
      15'b010_000011001011 : VALUE=19'b0000000_101100101101;
      15'b010_000011001100 : VALUE=19'b0000000_101100101101;
      15'b010_000011001101 : VALUE=19'b0000000_101100101101;
      15'b010_000011001110 : VALUE=19'b0000000_101100101101;
      15'b010_000011001111 : VALUE=19'b0000000_101100101100;
      15'b010_000011010000 : VALUE=19'b0000000_101100101100;
      15'b010_000011010001 : VALUE=19'b0000000_101100101100;
      15'b010_000011010010 : VALUE=19'b0000000_101100101100;
      15'b010_000011010011 : VALUE=19'b0000000_101100101100;
      15'b010_000011010100 : VALUE=19'b0000000_101100101100;
      15'b010_000011010101 : VALUE=19'b0000000_101100101011;
      15'b010_000011010110 : VALUE=19'b0000000_101100101011;
      15'b010_000011010111 : VALUE=19'b0000000_101100101011;
      15'b010_000011011000 : VALUE=19'b0000000_101100101011;
      15'b010_000011011001 : VALUE=19'b0000000_101100101011;
      15'b010_000011011010 : VALUE=19'b0000000_101100101011;
      15'b010_000011011011 : VALUE=19'b0000000_101100101010;
      15'b010_000011011100 : VALUE=19'b0000000_101100101010;
      15'b010_000011011101 : VALUE=19'b0000000_101100101010;
      15'b010_000011011110 : VALUE=19'b0000000_101100101010;
      15'b010_000011011111 : VALUE=19'b0000000_101100101010;
      15'b010_000011100000 : VALUE=19'b0000000_101100101010;
      15'b010_000011100001 : VALUE=19'b0000000_101100101001;
      15'b010_000011100010 : VALUE=19'b0000000_101100101001;
      15'b010_000011100011 : VALUE=19'b0000000_101100101001;
      15'b010_000011100100 : VALUE=19'b0000000_101100101001;
      15'b010_000011100101 : VALUE=19'b0000000_101100101001;
      15'b010_000011100110 : VALUE=19'b0000000_101100101000;
      15'b010_000011100111 : VALUE=19'b0000000_101100101000;
      15'b010_000011101000 : VALUE=19'b0000000_101100101000;
      15'b010_000011101001 : VALUE=19'b0000000_101100101000;
      15'b010_000011101010 : VALUE=19'b0000000_101100101000;
      15'b010_000011101011 : VALUE=19'b0000000_101100101000;
      15'b010_000011101100 : VALUE=19'b0000000_101100100111;
      15'b010_000011101101 : VALUE=19'b0000000_101100100111;
      15'b010_000011101110 : VALUE=19'b0000000_101100100111;
      15'b010_000011101111 : VALUE=19'b0000000_101100100111;
      15'b010_000011110000 : VALUE=19'b0000000_101100100111;
      15'b010_000011110001 : VALUE=19'b0000000_101100100111;
      15'b010_000011110010 : VALUE=19'b0000000_101100100110;
      15'b010_000011110011 : VALUE=19'b0000000_101100100110;
      15'b010_000011110100 : VALUE=19'b0000000_101100100110;
      15'b010_000011110101 : VALUE=19'b0000000_101100100110;
      15'b010_000011110110 : VALUE=19'b0000000_101100100110;
      15'b010_000011110111 : VALUE=19'b0000000_101100100110;
      15'b010_000011111000 : VALUE=19'b0000000_101100100101;
      15'b010_000011111001 : VALUE=19'b0000000_101100100101;
      15'b010_000011111010 : VALUE=19'b0000000_101100100101;
      15'b010_000011111011 : VALUE=19'b0000000_101100100101;
      15'b010_000011111100 : VALUE=19'b0000000_101100100101;
      15'b010_000011111101 : VALUE=19'b0000000_101100100101;
      15'b010_000011111110 : VALUE=19'b0000000_101100100100;
      15'b010_000011111111 : VALUE=19'b0000000_101100100100;
      15'b010_000100000000 : VALUE=19'b0000000_101100100100;
      15'b010_000100000001 : VALUE=19'b0000000_101100100100;
      15'b010_000100000010 : VALUE=19'b0000000_101100100100;
      15'b010_000100000011 : VALUE=19'b0000000_101100100100;
      15'b010_000100000100 : VALUE=19'b0000000_101100100011;
      15'b010_000100000101 : VALUE=19'b0000000_101100100011;
      15'b010_000100000110 : VALUE=19'b0000000_101100100011;
      15'b010_000100000111 : VALUE=19'b0000000_101100100011;
      15'b010_000100001000 : VALUE=19'b0000000_101100100011;
      15'b010_000100001001 : VALUE=19'b0000000_101100100011;
      15'b010_000100001010 : VALUE=19'b0000000_101100100010;
      15'b010_000100001011 : VALUE=19'b0000000_101100100010;
      15'b010_000100001100 : VALUE=19'b0000000_101100100010;
      15'b010_000100001101 : VALUE=19'b0000000_101100100010;
      15'b010_000100001110 : VALUE=19'b0000000_101100100010;
      15'b010_000100001111 : VALUE=19'b0000000_101100100010;
      15'b010_000100010000 : VALUE=19'b0000000_101100100001;
      15'b010_000100010001 : VALUE=19'b0000000_101100100001;
      15'b010_000100010010 : VALUE=19'b0000000_101100100001;
      15'b010_000100010011 : VALUE=19'b0000000_101100100001;
      15'b010_000100010100 : VALUE=19'b0000000_101100100001;
      15'b010_000100010101 : VALUE=19'b0000000_101100100001;
      15'b010_000100010110 : VALUE=19'b0000000_101100100000;
      15'b010_000100010111 : VALUE=19'b0000000_101100100000;
      15'b010_000100011000 : VALUE=19'b0000000_101100100000;
      15'b010_000100011001 : VALUE=19'b0000000_101100100000;
      15'b010_000100011010 : VALUE=19'b0000000_101100100000;
      15'b010_000100011011 : VALUE=19'b0000000_101100100000;
      15'b010_000100011100 : VALUE=19'b0000000_101100011111;
      15'b010_000100011101 : VALUE=19'b0000000_101100011111;
      15'b010_000100011110 : VALUE=19'b0000000_101100011111;
      15'b010_000100011111 : VALUE=19'b0000000_101100011111;
      15'b010_000100100000 : VALUE=19'b0000000_101100011111;
      15'b010_000100100001 : VALUE=19'b0000000_101100011111;
      15'b010_000100100010 : VALUE=19'b0000000_101100011110;
      15'b010_000100100011 : VALUE=19'b0000000_101100011110;
      15'b010_000100100100 : VALUE=19'b0000000_101100011110;
      15'b010_000100100101 : VALUE=19'b0000000_101100011110;
      15'b010_000100100110 : VALUE=19'b0000000_101100011110;
      15'b010_000100100111 : VALUE=19'b0000000_101100011110;
      15'b010_000100101000 : VALUE=19'b0000000_101100011101;
      15'b010_000100101001 : VALUE=19'b0000000_101100011101;
      15'b010_000100101010 : VALUE=19'b0000000_101100011101;
      15'b010_000100101011 : VALUE=19'b0000000_101100011101;
      15'b010_000100101100 : VALUE=19'b0000000_101100011101;
      15'b010_000100101101 : VALUE=19'b0000000_101100011101;
      15'b010_000100101110 : VALUE=19'b0000000_101100011100;
      15'b010_000100101111 : VALUE=19'b0000000_101100011100;
      15'b010_000100110000 : VALUE=19'b0000000_101100011100;
      15'b010_000100110001 : VALUE=19'b0000000_101100011100;
      15'b010_000100110010 : VALUE=19'b0000000_101100011100;
      15'b010_000100110011 : VALUE=19'b0000000_101100011100;
      15'b010_000100110100 : VALUE=19'b0000000_101100011011;
      15'b010_000100110101 : VALUE=19'b0000000_101100011011;
      15'b010_000100110110 : VALUE=19'b0000000_101100011011;
      15'b010_000100110111 : VALUE=19'b0000000_101100011011;
      15'b010_000100111000 : VALUE=19'b0000000_101100011011;
      15'b010_000100111001 : VALUE=19'b0000000_101100011011;
      15'b010_000100111010 : VALUE=19'b0000000_101100011010;
      15'b010_000100111011 : VALUE=19'b0000000_101100011010;
      15'b010_000100111100 : VALUE=19'b0000000_101100011010;
      15'b010_000100111101 : VALUE=19'b0000000_101100011010;
      15'b010_000100111110 : VALUE=19'b0000000_101100011010;
      15'b010_000100111111 : VALUE=19'b0000000_101100011010;
      15'b010_000101000000 : VALUE=19'b0000000_101100011001;
      15'b010_000101000001 : VALUE=19'b0000000_101100011001;
      15'b010_000101000010 : VALUE=19'b0000000_101100011001;
      15'b010_000101000011 : VALUE=19'b0000000_101100011001;
      15'b010_000101000100 : VALUE=19'b0000000_101100011001;
      15'b010_000101000101 : VALUE=19'b0000000_101100011001;
      15'b010_000101000110 : VALUE=19'b0000000_101100011000;
      15'b010_000101000111 : VALUE=19'b0000000_101100011000;
      15'b010_000101001000 : VALUE=19'b0000000_101100011000;
      15'b010_000101001001 : VALUE=19'b0000000_101100011000;
      15'b010_000101001010 : VALUE=19'b0000000_101100011000;
      15'b010_000101001011 : VALUE=19'b0000000_101100011000;
      15'b010_000101001100 : VALUE=19'b0000000_101100010111;
      15'b010_000101001101 : VALUE=19'b0000000_101100010111;
      15'b010_000101001110 : VALUE=19'b0000000_101100010111;
      15'b010_000101001111 : VALUE=19'b0000000_101100010111;
      15'b010_000101010000 : VALUE=19'b0000000_101100010111;
      15'b010_000101010001 : VALUE=19'b0000000_101100010111;
      15'b010_000101010010 : VALUE=19'b0000000_101100010110;
      15'b010_000101010011 : VALUE=19'b0000000_101100010110;
      15'b010_000101010100 : VALUE=19'b0000000_101100010110;
      15'b010_000101010101 : VALUE=19'b0000000_101100010110;
      15'b010_000101010110 : VALUE=19'b0000000_101100010110;
      15'b010_000101010111 : VALUE=19'b0000000_101100010110;
      15'b010_000101011000 : VALUE=19'b0000000_101100010101;
      15'b010_000101011001 : VALUE=19'b0000000_101100010101;
      15'b010_000101011010 : VALUE=19'b0000000_101100010101;
      15'b010_000101011011 : VALUE=19'b0000000_101100010101;
      15'b010_000101011100 : VALUE=19'b0000000_101100010101;
      15'b010_000101011101 : VALUE=19'b0000000_101100010101;
      15'b010_000101011110 : VALUE=19'b0000000_101100010100;
      15'b010_000101011111 : VALUE=19'b0000000_101100010100;
      15'b010_000101100000 : VALUE=19'b0000000_101100010100;
      15'b010_000101100001 : VALUE=19'b0000000_101100010100;
      15'b010_000101100010 : VALUE=19'b0000000_101100010100;
      15'b010_000101100011 : VALUE=19'b0000000_101100010100;
      15'b010_000101100100 : VALUE=19'b0000000_101100010011;
      15'b010_000101100101 : VALUE=19'b0000000_101100010011;
      15'b010_000101100110 : VALUE=19'b0000000_101100010011;
      15'b010_000101100111 : VALUE=19'b0000000_101100010011;
      15'b010_000101101000 : VALUE=19'b0000000_101100010011;
      15'b010_000101101001 : VALUE=19'b0000000_101100010011;
      15'b010_000101101010 : VALUE=19'b0000000_101100010010;
      15'b010_000101101011 : VALUE=19'b0000000_101100010010;
      15'b010_000101101100 : VALUE=19'b0000000_101100010010;
      15'b010_000101101101 : VALUE=19'b0000000_101100010010;
      15'b010_000101101110 : VALUE=19'b0000000_101100010010;
      15'b010_000101101111 : VALUE=19'b0000000_101100010010;
      15'b010_000101110000 : VALUE=19'b0000000_101100010001;
      15'b010_000101110001 : VALUE=19'b0000000_101100010001;
      15'b010_000101110010 : VALUE=19'b0000000_101100010001;
      15'b010_000101110011 : VALUE=19'b0000000_101100010001;
      15'b010_000101110100 : VALUE=19'b0000000_101100010001;
      15'b010_000101110101 : VALUE=19'b0000000_101100010001;
      15'b010_000101110110 : VALUE=19'b0000000_101100010000;
      15'b010_000101110111 : VALUE=19'b0000000_101100010000;
      15'b010_000101111000 : VALUE=19'b0000000_101100010000;
      15'b010_000101111001 : VALUE=19'b0000000_101100010000;
      15'b010_000101111010 : VALUE=19'b0000000_101100010000;
      15'b010_000101111011 : VALUE=19'b0000000_101100010000;
      15'b010_000101111100 : VALUE=19'b0000000_101100001111;
      15'b010_000101111101 : VALUE=19'b0000000_101100001111;
      15'b010_000101111110 : VALUE=19'b0000000_101100001111;
      15'b010_000101111111 : VALUE=19'b0000000_101100001111;
      15'b010_000110000000 : VALUE=19'b0000000_101100001111;
      15'b010_000110000001 : VALUE=19'b0000000_101100001111;
      15'b010_000110000010 : VALUE=19'b0000000_101100001110;
      15'b010_000110000011 : VALUE=19'b0000000_101100001110;
      15'b010_000110000100 : VALUE=19'b0000000_101100001110;
      15'b010_000110000101 : VALUE=19'b0000000_101100001110;
      15'b010_000110000110 : VALUE=19'b0000000_101100001110;
      15'b010_000110000111 : VALUE=19'b0000000_101100001110;
      15'b010_000110001000 : VALUE=19'b0000000_101100001101;
      15'b010_000110001001 : VALUE=19'b0000000_101100001101;
      15'b010_000110001010 : VALUE=19'b0000000_101100001101;
      15'b010_000110001011 : VALUE=19'b0000000_101100001101;
      15'b010_000110001100 : VALUE=19'b0000000_101100001101;
      15'b010_000110001101 : VALUE=19'b0000000_101100001101;
      15'b010_000110001110 : VALUE=19'b0000000_101100001100;
      15'b010_000110001111 : VALUE=19'b0000000_101100001100;
      15'b010_000110010000 : VALUE=19'b0000000_101100001100;
      15'b010_000110010001 : VALUE=19'b0000000_101100001100;
      15'b010_000110010010 : VALUE=19'b0000000_101100001100;
      15'b010_000110010011 : VALUE=19'b0000000_101100001100;
      15'b010_000110010100 : VALUE=19'b0000000_101100001011;
      15'b010_000110010101 : VALUE=19'b0000000_101100001011;
      15'b010_000110010110 : VALUE=19'b0000000_101100001011;
      15'b010_000110010111 : VALUE=19'b0000000_101100001011;
      15'b010_000110011000 : VALUE=19'b0000000_101100001011;
      15'b010_000110011001 : VALUE=19'b0000000_101100001011;
      15'b010_000110011010 : VALUE=19'b0000000_101100001010;
      15'b010_000110011011 : VALUE=19'b0000000_101100001010;
      15'b010_000110011100 : VALUE=19'b0000000_101100001010;
      15'b010_000110011101 : VALUE=19'b0000000_101100001010;
      15'b010_000110011110 : VALUE=19'b0000000_101100001010;
      15'b010_000110011111 : VALUE=19'b0000000_101100001010;
      15'b010_000110100000 : VALUE=19'b0000000_101100001001;
      15'b010_000110100001 : VALUE=19'b0000000_101100001001;
      15'b010_000110100010 : VALUE=19'b0000000_101100001001;
      15'b010_000110100011 : VALUE=19'b0000000_101100001001;
      15'b010_000110100100 : VALUE=19'b0000000_101100001001;
      15'b010_000110100101 : VALUE=19'b0000000_101100001001;
      15'b010_000110100110 : VALUE=19'b0000000_101100001000;
      15'b010_000110100111 : VALUE=19'b0000000_101100001000;
      15'b010_000110101000 : VALUE=19'b0000000_101100001000;
      15'b010_000110101001 : VALUE=19'b0000000_101100001000;
      15'b010_000110101010 : VALUE=19'b0000000_101100001000;
      15'b010_000110101011 : VALUE=19'b0000000_101100001000;
      15'b010_000110101100 : VALUE=19'b0000000_101100000111;
      15'b010_000110101101 : VALUE=19'b0000000_101100000111;
      15'b010_000110101110 : VALUE=19'b0000000_101100000111;
      15'b010_000110101111 : VALUE=19'b0000000_101100000111;
      15'b010_000110110000 : VALUE=19'b0000000_101100000111;
      15'b010_000110110001 : VALUE=19'b0000000_101100000111;
      15'b010_000110110010 : VALUE=19'b0000000_101100000111;
      15'b010_000110110011 : VALUE=19'b0000000_101100000110;
      15'b010_000110110100 : VALUE=19'b0000000_101100000110;
      15'b010_000110110101 : VALUE=19'b0000000_101100000110;
      15'b010_000110110110 : VALUE=19'b0000000_101100000110;
      15'b010_000110110111 : VALUE=19'b0000000_101100000110;
      15'b010_000110111000 : VALUE=19'b0000000_101100000110;
      15'b010_000110111001 : VALUE=19'b0000000_101100000101;
      15'b010_000110111010 : VALUE=19'b0000000_101100000101;
      15'b010_000110111011 : VALUE=19'b0000000_101100000101;
      15'b010_000110111100 : VALUE=19'b0000000_101100000101;
      15'b010_000110111101 : VALUE=19'b0000000_101100000101;
      15'b010_000110111110 : VALUE=19'b0000000_101100000101;
      15'b010_000110111111 : VALUE=19'b0000000_101100000100;
      15'b010_000111000000 : VALUE=19'b0000000_101100000100;
      15'b010_000111000001 : VALUE=19'b0000000_101100000100;
      15'b010_000111000010 : VALUE=19'b0000000_101100000100;
      15'b010_000111000011 : VALUE=19'b0000000_101100000100;
      15'b010_000111000100 : VALUE=19'b0000000_101100000100;
      15'b010_000111000101 : VALUE=19'b0000000_101100000011;
      15'b010_000111000110 : VALUE=19'b0000000_101100000011;
      15'b010_000111000111 : VALUE=19'b0000000_101100000011;
      15'b010_000111001000 : VALUE=19'b0000000_101100000011;
      15'b010_000111001001 : VALUE=19'b0000000_101100000011;
      15'b010_000111001010 : VALUE=19'b0000000_101100000011;
      15'b010_000111001011 : VALUE=19'b0000000_101100000010;
      15'b010_000111001100 : VALUE=19'b0000000_101100000010;
      15'b010_000111001101 : VALUE=19'b0000000_101100000010;
      15'b010_000111001110 : VALUE=19'b0000000_101100000010;
      15'b010_000111001111 : VALUE=19'b0000000_101100000010;
      15'b010_000111010000 : VALUE=19'b0000000_101100000010;
      15'b010_000111010001 : VALUE=19'b0000000_101100000001;
      15'b010_000111010010 : VALUE=19'b0000000_101100000001;
      15'b010_000111010011 : VALUE=19'b0000000_101100000001;
      15'b010_000111010100 : VALUE=19'b0000000_101100000001;
      15'b010_000111010101 : VALUE=19'b0000000_101100000001;
      15'b010_000111010110 : VALUE=19'b0000000_101100000001;
      15'b010_000111010111 : VALUE=19'b0000000_101100000000;
      15'b010_000111011000 : VALUE=19'b0000000_101100000000;
      15'b010_000111011001 : VALUE=19'b0000000_101100000000;
      15'b010_000111011010 : VALUE=19'b0000000_101100000000;
      15'b010_000111011011 : VALUE=19'b0000000_101100000000;
      15'b010_000111011100 : VALUE=19'b0000000_101100000000;
      15'b010_000111011101 : VALUE=19'b0000000_101011111111;
      15'b010_000111011110 : VALUE=19'b0000000_101011111111;
      15'b010_000111011111 : VALUE=19'b0000000_101011111111;
      15'b010_000111100000 : VALUE=19'b0000000_101011111111;
      15'b010_000111100001 : VALUE=19'b0000000_101011111111;
      15'b010_000111100010 : VALUE=19'b0000000_101011111111;
      15'b010_000111100011 : VALUE=19'b0000000_101011111111;
      15'b010_000111100100 : VALUE=19'b0000000_101011111110;
      15'b010_000111100101 : VALUE=19'b0000000_101011111110;
      15'b010_000111100110 : VALUE=19'b0000000_101011111110;
      15'b010_000111100111 : VALUE=19'b0000000_101011111110;
      15'b010_000111101000 : VALUE=19'b0000000_101011111110;
      15'b010_000111101001 : VALUE=19'b0000000_101011111110;
      15'b010_000111101010 : VALUE=19'b0000000_101011111101;
      15'b010_000111101011 : VALUE=19'b0000000_101011111101;
      15'b010_000111101100 : VALUE=19'b0000000_101011111101;
      15'b010_000111101101 : VALUE=19'b0000000_101011111101;
      15'b010_000111101110 : VALUE=19'b0000000_101011111101;
      15'b010_000111101111 : VALUE=19'b0000000_101011111101;
      15'b010_000111110000 : VALUE=19'b0000000_101011111100;
      15'b010_000111110001 : VALUE=19'b0000000_101011111100;
      15'b010_000111110010 : VALUE=19'b0000000_101011111100;
      15'b010_000111110011 : VALUE=19'b0000000_101011111100;
      15'b010_000111110100 : VALUE=19'b0000000_101011111100;
      15'b010_000111110101 : VALUE=19'b0000000_101011111100;
      15'b010_000111110110 : VALUE=19'b0000000_101011111011;
      15'b010_000111110111 : VALUE=19'b0000000_101011111011;
      15'b010_000111111000 : VALUE=19'b0000000_101011111011;
      15'b010_000111111001 : VALUE=19'b0000000_101011111011;
      15'b010_000111111010 : VALUE=19'b0000000_101011111011;
      15'b010_000111111011 : VALUE=19'b0000000_101011111011;
      15'b010_000111111100 : VALUE=19'b0000000_101011111010;
      15'b010_000111111101 : VALUE=19'b0000000_101011111010;
      15'b010_000111111110 : VALUE=19'b0000000_101011111010;
      15'b010_000111111111 : VALUE=19'b0000000_101011111010;
      15'b010_001000000000 : VALUE=19'b0000000_101011111010;
      15'b010_001000000001 : VALUE=19'b0000000_101011111010;
      15'b010_001000000010 : VALUE=19'b0000000_101011111010;
      15'b010_001000000011 : VALUE=19'b0000000_101011111001;
      15'b010_001000000100 : VALUE=19'b0000000_101011111001;
      15'b010_001000000101 : VALUE=19'b0000000_101011111001;
      15'b010_001000000110 : VALUE=19'b0000000_101011111001;
      15'b010_001000000111 : VALUE=19'b0000000_101011111001;
      15'b010_001000001000 : VALUE=19'b0000000_101011111001;
      15'b010_001000001001 : VALUE=19'b0000000_101011111000;
      15'b010_001000001010 : VALUE=19'b0000000_101011111000;
      15'b010_001000001011 : VALUE=19'b0000000_101011111000;
      15'b010_001000001100 : VALUE=19'b0000000_101011111000;
      15'b010_001000001101 : VALUE=19'b0000000_101011111000;
      15'b010_001000001110 : VALUE=19'b0000000_101011111000;
      15'b010_001000001111 : VALUE=19'b0000000_101011110111;
      15'b010_001000010000 : VALUE=19'b0000000_101011110111;
      15'b010_001000010001 : VALUE=19'b0000000_101011110111;
      15'b010_001000010010 : VALUE=19'b0000000_101011110111;
      15'b010_001000010011 : VALUE=19'b0000000_101011110111;
      15'b010_001000010100 : VALUE=19'b0000000_101011110111;
      15'b010_001000010101 : VALUE=19'b0000000_101011110110;
      15'b010_001000010110 : VALUE=19'b0000000_101011110110;
      15'b010_001000010111 : VALUE=19'b0000000_101011110110;
      15'b010_001000011000 : VALUE=19'b0000000_101011110110;
      15'b010_001000011001 : VALUE=19'b0000000_101011110110;
      15'b010_001000011010 : VALUE=19'b0000000_101011110110;
      15'b010_001000011011 : VALUE=19'b0000000_101011110101;
      15'b010_001000011100 : VALUE=19'b0000000_101011110101;
      15'b010_001000011101 : VALUE=19'b0000000_101011110101;
      15'b010_001000011110 : VALUE=19'b0000000_101011110101;
      15'b010_001000011111 : VALUE=19'b0000000_101011110101;
      15'b010_001000100000 : VALUE=19'b0000000_101011110101;
      15'b010_001000100001 : VALUE=19'b0000000_101011110101;
      15'b010_001000100010 : VALUE=19'b0000000_101011110100;
      15'b010_001000100011 : VALUE=19'b0000000_101011110100;
      15'b010_001000100100 : VALUE=19'b0000000_101011110100;
      15'b010_001000100101 : VALUE=19'b0000000_101011110100;
      15'b010_001000100110 : VALUE=19'b0000000_101011110100;
      15'b010_001000100111 : VALUE=19'b0000000_101011110100;
      15'b010_001000101000 : VALUE=19'b0000000_101011110011;
      15'b010_001000101001 : VALUE=19'b0000000_101011110011;
      15'b010_001000101010 : VALUE=19'b0000000_101011110011;
      15'b010_001000101011 : VALUE=19'b0000000_101011110011;
      15'b010_001000101100 : VALUE=19'b0000000_101011110011;
      15'b010_001000101101 : VALUE=19'b0000000_101011110011;
      15'b010_001000101110 : VALUE=19'b0000000_101011110010;
      15'b010_001000101111 : VALUE=19'b0000000_101011110010;
      15'b010_001000110000 : VALUE=19'b0000000_101011110010;
      15'b010_001000110001 : VALUE=19'b0000000_101011110010;
      15'b010_001000110010 : VALUE=19'b0000000_101011110010;
      15'b010_001000110011 : VALUE=19'b0000000_101011110010;
      15'b010_001000110100 : VALUE=19'b0000000_101011110001;
      15'b010_001000110101 : VALUE=19'b0000000_101011110001;
      15'b010_001000110110 : VALUE=19'b0000000_101011110001;
      15'b010_001000110111 : VALUE=19'b0000000_101011110001;
      15'b010_001000111000 : VALUE=19'b0000000_101011110001;
      15'b010_001000111001 : VALUE=19'b0000000_101011110001;
      15'b010_001000111010 : VALUE=19'b0000000_101011110001;
      15'b010_001000111011 : VALUE=19'b0000000_101011110000;
      15'b010_001000111100 : VALUE=19'b0000000_101011110000;
      15'b010_001000111101 : VALUE=19'b0000000_101011110000;
      15'b010_001000111110 : VALUE=19'b0000000_101011110000;
      15'b010_001000111111 : VALUE=19'b0000000_101011110000;
      15'b010_001001000000 : VALUE=19'b0000000_101011110000;
      15'b010_001001000001 : VALUE=19'b0000000_101011101111;
      15'b010_001001000010 : VALUE=19'b0000000_101011101111;
      15'b010_001001000011 : VALUE=19'b0000000_101011101111;
      15'b010_001001000100 : VALUE=19'b0000000_101011101111;
      15'b010_001001000101 : VALUE=19'b0000000_101011101111;
      15'b010_001001000110 : VALUE=19'b0000000_101011101111;
      15'b010_001001000111 : VALUE=19'b0000000_101011101110;
      15'b010_001001001000 : VALUE=19'b0000000_101011101110;
      15'b010_001001001001 : VALUE=19'b0000000_101011101110;
      15'b010_001001001010 : VALUE=19'b0000000_101011101110;
      15'b010_001001001011 : VALUE=19'b0000000_101011101110;
      15'b010_001001001100 : VALUE=19'b0000000_101011101110;
      15'b010_001001001101 : VALUE=19'b0000000_101011101101;
      15'b010_001001001110 : VALUE=19'b0000000_101011101101;
      15'b010_001001001111 : VALUE=19'b0000000_101011101101;
      15'b010_001001010000 : VALUE=19'b0000000_101011101101;
      15'b010_001001010001 : VALUE=19'b0000000_101011101101;
      15'b010_001001010010 : VALUE=19'b0000000_101011101101;
      15'b010_001001010011 : VALUE=19'b0000000_101011101101;
      15'b010_001001010100 : VALUE=19'b0000000_101011101100;
      15'b010_001001010101 : VALUE=19'b0000000_101011101100;
      15'b010_001001010110 : VALUE=19'b0000000_101011101100;
      15'b010_001001010111 : VALUE=19'b0000000_101011101100;
      15'b010_001001011000 : VALUE=19'b0000000_101011101100;
      15'b010_001001011001 : VALUE=19'b0000000_101011101100;
      15'b010_001001011010 : VALUE=19'b0000000_101011101011;
      15'b010_001001011011 : VALUE=19'b0000000_101011101011;
      15'b010_001001011100 : VALUE=19'b0000000_101011101011;
      15'b010_001001011101 : VALUE=19'b0000000_101011101011;
      15'b010_001001011110 : VALUE=19'b0000000_101011101011;
      15'b010_001001011111 : VALUE=19'b0000000_101011101011;
      15'b010_001001100000 : VALUE=19'b0000000_101011101010;
      15'b010_001001100001 : VALUE=19'b0000000_101011101010;
      15'b010_001001100010 : VALUE=19'b0000000_101011101010;
      15'b010_001001100011 : VALUE=19'b0000000_101011101010;
      15'b010_001001100100 : VALUE=19'b0000000_101011101010;
      15'b010_001001100101 : VALUE=19'b0000000_101011101010;
      15'b010_001001100110 : VALUE=19'b0000000_101011101010;
      15'b010_001001100111 : VALUE=19'b0000000_101011101001;
      15'b010_001001101000 : VALUE=19'b0000000_101011101001;
      15'b010_001001101001 : VALUE=19'b0000000_101011101001;
      15'b010_001001101010 : VALUE=19'b0000000_101011101001;
      15'b010_001001101011 : VALUE=19'b0000000_101011101001;
      15'b010_001001101100 : VALUE=19'b0000000_101011101001;
      15'b010_001001101101 : VALUE=19'b0000000_101011101000;
      15'b010_001001101110 : VALUE=19'b0000000_101011101000;
      15'b010_001001101111 : VALUE=19'b0000000_101011101000;
      15'b010_001001110000 : VALUE=19'b0000000_101011101000;
      15'b010_001001110001 : VALUE=19'b0000000_101011101000;
      15'b010_001001110010 : VALUE=19'b0000000_101011101000;
      15'b010_001001110011 : VALUE=19'b0000000_101011100111;
      15'b010_001001110100 : VALUE=19'b0000000_101011100111;
      15'b010_001001110101 : VALUE=19'b0000000_101011100111;
      15'b010_001001110110 : VALUE=19'b0000000_101011100111;
      15'b010_001001110111 : VALUE=19'b0000000_101011100111;
      15'b010_001001111000 : VALUE=19'b0000000_101011100111;
      15'b010_001001111001 : VALUE=19'b0000000_101011100111;
      15'b010_001001111010 : VALUE=19'b0000000_101011100110;
      15'b010_001001111011 : VALUE=19'b0000000_101011100110;
      15'b010_001001111100 : VALUE=19'b0000000_101011100110;
      15'b010_001001111101 : VALUE=19'b0000000_101011100110;
      15'b010_001001111110 : VALUE=19'b0000000_101011100110;
      15'b010_001001111111 : VALUE=19'b0000000_101011100110;
      15'b010_001010000000 : VALUE=19'b0000000_101011100101;
      15'b010_001010000001 : VALUE=19'b0000000_101011100101;
      15'b010_001010000010 : VALUE=19'b0000000_101011100101;
      15'b010_001010000011 : VALUE=19'b0000000_101011100101;
      15'b010_001010000100 : VALUE=19'b0000000_101011100101;
      15'b010_001010000101 : VALUE=19'b0000000_101011100101;
      15'b010_001010000110 : VALUE=19'b0000000_101011100100;
      15'b010_001010000111 : VALUE=19'b0000000_101011100100;
      15'b010_001010001000 : VALUE=19'b0000000_101011100100;
      15'b010_001010001001 : VALUE=19'b0000000_101011100100;
      15'b010_001010001010 : VALUE=19'b0000000_101011100100;
      15'b010_001010001011 : VALUE=19'b0000000_101011100100;
      15'b010_001010001100 : VALUE=19'b0000000_101011100100;
      15'b010_001010001101 : VALUE=19'b0000000_101011100011;
      15'b010_001010001110 : VALUE=19'b0000000_101011100011;
      15'b010_001010001111 : VALUE=19'b0000000_101011100011;
      15'b010_001010010000 : VALUE=19'b0000000_101011100011;
      15'b010_001010010001 : VALUE=19'b0000000_101011100011;
      15'b010_001010010010 : VALUE=19'b0000000_101011100011;
      15'b010_001010010011 : VALUE=19'b0000000_101011100010;
      15'b010_001010010100 : VALUE=19'b0000000_101011100010;
      15'b010_001010010101 : VALUE=19'b0000000_101011100010;
      15'b010_001010010110 : VALUE=19'b0000000_101011100010;
      15'b010_001010010111 : VALUE=19'b0000000_101011100010;
      15'b010_001010011000 : VALUE=19'b0000000_101011100010;
      15'b010_001010011001 : VALUE=19'b0000000_101011100001;
      15'b010_001010011010 : VALUE=19'b0000000_101011100001;
      15'b010_001010011011 : VALUE=19'b0000000_101011100001;
      15'b010_001010011100 : VALUE=19'b0000000_101011100001;
      15'b010_001010011101 : VALUE=19'b0000000_101011100001;
      15'b010_001010011110 : VALUE=19'b0000000_101011100001;
      15'b010_001010011111 : VALUE=19'b0000000_101011100001;
      15'b010_001010100000 : VALUE=19'b0000000_101011100000;
      15'b010_001010100001 : VALUE=19'b0000000_101011100000;
      15'b010_001010100010 : VALUE=19'b0000000_101011100000;
      15'b010_001010100011 : VALUE=19'b0000000_101011100000;
      15'b010_001010100100 : VALUE=19'b0000000_101011100000;
      15'b010_001010100101 : VALUE=19'b0000000_101011100000;
      15'b010_001010100110 : VALUE=19'b0000000_101011011111;
      15'b010_001010100111 : VALUE=19'b0000000_101011011111;
      15'b010_001010101000 : VALUE=19'b0000000_101011011111;
      15'b010_001010101001 : VALUE=19'b0000000_101011011111;
      15'b010_001010101010 : VALUE=19'b0000000_101011011111;
      15'b010_001010101011 : VALUE=19'b0000000_101011011111;
      15'b010_001010101100 : VALUE=19'b0000000_101011011110;
      15'b010_001010101101 : VALUE=19'b0000000_101011011110;
      15'b010_001010101110 : VALUE=19'b0000000_101011011110;
      15'b010_001010101111 : VALUE=19'b0000000_101011011110;
      15'b010_001010110000 : VALUE=19'b0000000_101011011110;
      15'b010_001010110001 : VALUE=19'b0000000_101011011110;
      15'b010_001010110010 : VALUE=19'b0000000_101011011110;
      15'b010_001010110011 : VALUE=19'b0000000_101011011101;
      15'b010_001010110100 : VALUE=19'b0000000_101011011101;
      15'b010_001010110101 : VALUE=19'b0000000_101011011101;
      15'b010_001010110110 : VALUE=19'b0000000_101011011101;
      15'b010_001010110111 : VALUE=19'b0000000_101011011101;
      15'b010_001010111000 : VALUE=19'b0000000_101011011101;
      15'b010_001010111001 : VALUE=19'b0000000_101011011100;
      15'b010_001010111010 : VALUE=19'b0000000_101011011100;
      15'b010_001010111011 : VALUE=19'b0000000_101011011100;
      15'b010_001010111100 : VALUE=19'b0000000_101011011100;
      15'b010_001010111101 : VALUE=19'b0000000_101011011100;
      15'b010_001010111110 : VALUE=19'b0000000_101011011100;
      15'b010_001010111111 : VALUE=19'b0000000_101011011100;
      15'b010_001011000000 : VALUE=19'b0000000_101011011011;
      15'b010_001011000001 : VALUE=19'b0000000_101011011011;
      15'b010_001011000010 : VALUE=19'b0000000_101011011011;
      15'b010_001011000011 : VALUE=19'b0000000_101011011011;
      15'b010_001011000100 : VALUE=19'b0000000_101011011011;
      15'b010_001011000101 : VALUE=19'b0000000_101011011011;
      15'b010_001011000110 : VALUE=19'b0000000_101011011010;
      15'b010_001011000111 : VALUE=19'b0000000_101011011010;
      15'b010_001011001000 : VALUE=19'b0000000_101011011010;
      15'b010_001011001001 : VALUE=19'b0000000_101011011010;
      15'b010_001011001010 : VALUE=19'b0000000_101011011010;
      15'b010_001011001011 : VALUE=19'b0000000_101011011010;
      15'b010_001011001100 : VALUE=19'b0000000_101011011001;
      15'b010_001011001101 : VALUE=19'b0000000_101011011001;
      15'b010_001011001110 : VALUE=19'b0000000_101011011001;
      15'b010_001011001111 : VALUE=19'b0000000_101011011001;
      15'b010_001011010000 : VALUE=19'b0000000_101011011001;
      15'b010_001011010001 : VALUE=19'b0000000_101011011001;
      15'b010_001011010010 : VALUE=19'b0000000_101011011001;
      15'b010_001011010011 : VALUE=19'b0000000_101011011000;
      15'b010_001011010100 : VALUE=19'b0000000_101011011000;
      15'b010_001011010101 : VALUE=19'b0000000_101011011000;
      15'b010_001011010110 : VALUE=19'b0000000_101011011000;
      15'b010_001011010111 : VALUE=19'b0000000_101011011000;
      15'b010_001011011000 : VALUE=19'b0000000_101011011000;
      15'b010_001011011001 : VALUE=19'b0000000_101011010111;
      15'b010_001011011010 : VALUE=19'b0000000_101011010111;
      15'b010_001011011011 : VALUE=19'b0000000_101011010111;
      15'b010_001011011100 : VALUE=19'b0000000_101011010111;
      15'b010_001011011101 : VALUE=19'b0000000_101011010111;
      15'b010_001011011110 : VALUE=19'b0000000_101011010111;
      15'b010_001011011111 : VALUE=19'b0000000_101011010111;
      15'b010_001011100000 : VALUE=19'b0000000_101011010110;
      15'b010_001011100001 : VALUE=19'b0000000_101011010110;
      15'b010_001011100010 : VALUE=19'b0000000_101011010110;
      15'b010_001011100011 : VALUE=19'b0000000_101011010110;
      15'b010_001011100100 : VALUE=19'b0000000_101011010110;
      15'b010_001011100101 : VALUE=19'b0000000_101011010110;
      15'b010_001011100110 : VALUE=19'b0000000_101011010101;
      15'b010_001011100111 : VALUE=19'b0000000_101011010101;
      15'b010_001011101000 : VALUE=19'b0000000_101011010101;
      15'b010_001011101001 : VALUE=19'b0000000_101011010101;
      15'b010_001011101010 : VALUE=19'b0000000_101011010101;
      15'b010_001011101011 : VALUE=19'b0000000_101011010101;
      15'b010_001011101100 : VALUE=19'b0000000_101011010100;
      15'b010_001011101101 : VALUE=19'b0000000_101011010100;
      15'b010_001011101110 : VALUE=19'b0000000_101011010100;
      15'b010_001011101111 : VALUE=19'b0000000_101011010100;
      15'b010_001011110000 : VALUE=19'b0000000_101011010100;
      15'b010_001011110001 : VALUE=19'b0000000_101011010100;
      15'b010_001011110010 : VALUE=19'b0000000_101011010100;
      15'b010_001011110011 : VALUE=19'b0000000_101011010011;
      15'b010_001011110100 : VALUE=19'b0000000_101011010011;
      15'b010_001011110101 : VALUE=19'b0000000_101011010011;
      15'b010_001011110110 : VALUE=19'b0000000_101011010011;
      15'b010_001011110111 : VALUE=19'b0000000_101011010011;
      15'b010_001011111000 : VALUE=19'b0000000_101011010011;
      15'b010_001011111001 : VALUE=19'b0000000_101011010010;
      15'b010_001011111010 : VALUE=19'b0000000_101011010010;
      15'b010_001011111011 : VALUE=19'b0000000_101011010010;
      15'b010_001011111100 : VALUE=19'b0000000_101011010010;
      15'b010_001011111101 : VALUE=19'b0000000_101011010010;
      15'b010_001011111110 : VALUE=19'b0000000_101011010010;
      15'b010_001011111111 : VALUE=19'b0000000_101011010010;
      15'b010_001100000000 : VALUE=19'b0000000_101011010001;
      15'b010_001100000001 : VALUE=19'b0000000_101011010001;
      15'b010_001100000010 : VALUE=19'b0000000_101011010001;
      15'b010_001100000011 : VALUE=19'b0000000_101011010001;
      15'b010_001100000100 : VALUE=19'b0000000_101011010001;
      15'b010_001100000101 : VALUE=19'b0000000_101011010001;
      15'b010_001100000110 : VALUE=19'b0000000_101011010000;
      15'b010_001100000111 : VALUE=19'b0000000_101011010000;
      15'b010_001100001000 : VALUE=19'b0000000_101011010000;
      15'b010_001100001001 : VALUE=19'b0000000_101011010000;
      15'b010_001100001010 : VALUE=19'b0000000_101011010000;
      15'b010_001100001011 : VALUE=19'b0000000_101011010000;
      15'b010_001100001100 : VALUE=19'b0000000_101011010000;
      15'b010_001100001101 : VALUE=19'b0000000_101011001111;
      15'b010_001100001110 : VALUE=19'b0000000_101011001111;
      15'b010_001100001111 : VALUE=19'b0000000_101011001111;
      15'b010_001100010000 : VALUE=19'b0000000_101011001111;
      15'b010_001100010001 : VALUE=19'b0000000_101011001111;
      15'b010_001100010010 : VALUE=19'b0000000_101011001111;
      15'b010_001100010011 : VALUE=19'b0000000_101011001110;
      15'b010_001100010100 : VALUE=19'b0000000_101011001110;
      15'b010_001100010101 : VALUE=19'b0000000_101011001110;
      15'b010_001100010110 : VALUE=19'b0000000_101011001110;
      15'b010_001100010111 : VALUE=19'b0000000_101011001110;
      15'b010_001100011000 : VALUE=19'b0000000_101011001110;
      15'b010_001100011001 : VALUE=19'b0000000_101011001110;
      15'b010_001100011010 : VALUE=19'b0000000_101011001101;
      15'b010_001100011011 : VALUE=19'b0000000_101011001101;
      15'b010_001100011100 : VALUE=19'b0000000_101011001101;
      15'b010_001100011101 : VALUE=19'b0000000_101011001101;
      15'b010_001100011110 : VALUE=19'b0000000_101011001101;
      15'b010_001100011111 : VALUE=19'b0000000_101011001101;
      15'b010_001100100000 : VALUE=19'b0000000_101011001100;
      15'b010_001100100001 : VALUE=19'b0000000_101011001100;
      15'b010_001100100010 : VALUE=19'b0000000_101011001100;
      15'b010_001100100011 : VALUE=19'b0000000_101011001100;
      15'b010_001100100100 : VALUE=19'b0000000_101011001100;
      15'b010_001100100101 : VALUE=19'b0000000_101011001100;
      15'b010_001100100110 : VALUE=19'b0000000_101011001100;
      15'b010_001100100111 : VALUE=19'b0000000_101011001011;
      15'b010_001100101000 : VALUE=19'b0000000_101011001011;
      15'b010_001100101001 : VALUE=19'b0000000_101011001011;
      15'b010_001100101010 : VALUE=19'b0000000_101011001011;
      15'b010_001100101011 : VALUE=19'b0000000_101011001011;
      15'b010_001100101100 : VALUE=19'b0000000_101011001011;
      15'b010_001100101101 : VALUE=19'b0000000_101011001010;
      15'b010_001100101110 : VALUE=19'b0000000_101011001010;
      15'b010_001100101111 : VALUE=19'b0000000_101011001010;
      15'b010_001100110000 : VALUE=19'b0000000_101011001010;
      15'b010_001100110001 : VALUE=19'b0000000_101011001010;
      15'b010_001100110010 : VALUE=19'b0000000_101011001010;
      15'b010_001100110011 : VALUE=19'b0000000_101011001010;
      15'b010_001100110100 : VALUE=19'b0000000_101011001001;
      15'b010_001100110101 : VALUE=19'b0000000_101011001001;
      15'b010_001100110110 : VALUE=19'b0000000_101011001001;
      15'b010_001100110111 : VALUE=19'b0000000_101011001001;
      15'b010_001100111000 : VALUE=19'b0000000_101011001001;
      15'b010_001100111001 : VALUE=19'b0000000_101011001001;
      15'b010_001100111010 : VALUE=19'b0000000_101011001000;
      15'b010_001100111011 : VALUE=19'b0000000_101011001000;
      15'b010_001100111100 : VALUE=19'b0000000_101011001000;
      15'b010_001100111101 : VALUE=19'b0000000_101011001000;
      15'b010_001100111110 : VALUE=19'b0000000_101011001000;
      15'b010_001100111111 : VALUE=19'b0000000_101011001000;
      15'b010_001101000000 : VALUE=19'b0000000_101011001000;
      15'b010_001101000001 : VALUE=19'b0000000_101011000111;
      15'b010_001101000010 : VALUE=19'b0000000_101011000111;
      15'b010_001101000011 : VALUE=19'b0000000_101011000111;
      15'b010_001101000100 : VALUE=19'b0000000_101011000111;
      15'b010_001101000101 : VALUE=19'b0000000_101011000111;
      15'b010_001101000110 : VALUE=19'b0000000_101011000111;
      15'b010_001101000111 : VALUE=19'b0000000_101011000110;
      15'b010_001101001000 : VALUE=19'b0000000_101011000110;
      15'b010_001101001001 : VALUE=19'b0000000_101011000110;
      15'b010_001101001010 : VALUE=19'b0000000_101011000110;
      15'b010_001101001011 : VALUE=19'b0000000_101011000110;
      15'b010_001101001100 : VALUE=19'b0000000_101011000110;
      15'b010_001101001101 : VALUE=19'b0000000_101011000110;
      15'b010_001101001110 : VALUE=19'b0000000_101011000101;
      15'b010_001101001111 : VALUE=19'b0000000_101011000101;
      15'b010_001101010000 : VALUE=19'b0000000_101011000101;
      15'b010_001101010001 : VALUE=19'b0000000_101011000101;
      15'b010_001101010010 : VALUE=19'b0000000_101011000101;
      15'b010_001101010011 : VALUE=19'b0000000_101011000101;
      15'b010_001101010100 : VALUE=19'b0000000_101011000101;
      15'b010_001101010101 : VALUE=19'b0000000_101011000100;
      15'b010_001101010110 : VALUE=19'b0000000_101011000100;
      15'b010_001101010111 : VALUE=19'b0000000_101011000100;
      15'b010_001101011000 : VALUE=19'b0000000_101011000100;
      15'b010_001101011001 : VALUE=19'b0000000_101011000100;
      15'b010_001101011010 : VALUE=19'b0000000_101011000100;
      15'b010_001101011011 : VALUE=19'b0000000_101011000011;
      15'b010_001101011100 : VALUE=19'b0000000_101011000011;
      15'b010_001101011101 : VALUE=19'b0000000_101011000011;
      15'b010_001101011110 : VALUE=19'b0000000_101011000011;
      15'b010_001101011111 : VALUE=19'b0000000_101011000011;
      15'b010_001101100000 : VALUE=19'b0000000_101011000011;
      15'b010_001101100001 : VALUE=19'b0000000_101011000011;
      15'b010_001101100010 : VALUE=19'b0000000_101011000010;
      15'b010_001101100011 : VALUE=19'b0000000_101011000010;
      15'b010_001101100100 : VALUE=19'b0000000_101011000010;
      15'b010_001101100101 : VALUE=19'b0000000_101011000010;
      15'b010_001101100110 : VALUE=19'b0000000_101011000010;
      15'b010_001101100111 : VALUE=19'b0000000_101011000010;
      15'b010_001101101000 : VALUE=19'b0000000_101011000001;
      15'b010_001101101001 : VALUE=19'b0000000_101011000001;
      15'b010_001101101010 : VALUE=19'b0000000_101011000001;
      15'b010_001101101011 : VALUE=19'b0000000_101011000001;
      15'b010_001101101100 : VALUE=19'b0000000_101011000001;
      15'b010_001101101101 : VALUE=19'b0000000_101011000001;
      15'b010_001101101110 : VALUE=19'b0000000_101011000001;
      15'b010_001101101111 : VALUE=19'b0000000_101011000000;
      15'b010_001101110000 : VALUE=19'b0000000_101011000000;
      15'b010_001101110001 : VALUE=19'b0000000_101011000000;
      15'b010_001101110010 : VALUE=19'b0000000_101011000000;
      15'b010_001101110011 : VALUE=19'b0000000_101011000000;
      15'b010_001101110100 : VALUE=19'b0000000_101011000000;
      15'b010_001101110101 : VALUE=19'b0000000_101010111111;
      15'b010_001101110110 : VALUE=19'b0000000_101010111111;
      15'b010_001101110111 : VALUE=19'b0000000_101010111111;
      15'b010_001101111000 : VALUE=19'b0000000_101010111111;
      15'b010_001101111001 : VALUE=19'b0000000_101010111111;
      15'b010_001101111010 : VALUE=19'b0000000_101010111111;
      15'b010_001101111011 : VALUE=19'b0000000_101010111111;
      15'b010_001101111100 : VALUE=19'b0000000_101010111110;
      15'b010_001101111101 : VALUE=19'b0000000_101010111110;
      15'b010_001101111110 : VALUE=19'b0000000_101010111110;
      15'b010_001101111111 : VALUE=19'b0000000_101010111110;
      15'b010_001110000000 : VALUE=19'b0000000_101010111110;
      15'b010_001110000001 : VALUE=19'b0000000_101010111110;
      15'b010_001110000010 : VALUE=19'b0000000_101010111110;
      15'b010_001110000011 : VALUE=19'b0000000_101010111101;
      15'b010_001110000100 : VALUE=19'b0000000_101010111101;
      15'b010_001110000101 : VALUE=19'b0000000_101010111101;
      15'b010_001110000110 : VALUE=19'b0000000_101010111101;
      15'b010_001110000111 : VALUE=19'b0000000_101010111101;
      15'b010_001110001000 : VALUE=19'b0000000_101010111101;
      15'b010_001110001001 : VALUE=19'b0000000_101010111100;
      15'b010_001110001010 : VALUE=19'b0000000_101010111100;
      15'b010_001110001011 : VALUE=19'b0000000_101010111100;
      15'b010_001110001100 : VALUE=19'b0000000_101010111100;
      15'b010_001110001101 : VALUE=19'b0000000_101010111100;
      15'b010_001110001110 : VALUE=19'b0000000_101010111100;
      15'b010_001110001111 : VALUE=19'b0000000_101010111100;
      15'b010_001110010000 : VALUE=19'b0000000_101010111011;
      15'b010_001110010001 : VALUE=19'b0000000_101010111011;
      15'b010_001110010010 : VALUE=19'b0000000_101010111011;
      15'b010_001110010011 : VALUE=19'b0000000_101010111011;
      15'b010_001110010100 : VALUE=19'b0000000_101010111011;
      15'b010_001110010101 : VALUE=19'b0000000_101010111011;
      15'b010_001110010110 : VALUE=19'b0000000_101010111011;
      15'b010_001110010111 : VALUE=19'b0000000_101010111010;
      15'b010_001110011000 : VALUE=19'b0000000_101010111010;
      15'b010_001110011001 : VALUE=19'b0000000_101010111010;
      15'b010_001110011010 : VALUE=19'b0000000_101010111010;
      15'b010_001110011011 : VALUE=19'b0000000_101010111010;
      15'b010_001110011100 : VALUE=19'b0000000_101010111010;
      15'b010_001110011101 : VALUE=19'b0000000_101010111001;
      15'b010_001110011110 : VALUE=19'b0000000_101010111001;
      15'b010_001110011111 : VALUE=19'b0000000_101010111001;
      15'b010_001110100000 : VALUE=19'b0000000_101010111001;
      15'b010_001110100001 : VALUE=19'b0000000_101010111001;
      15'b010_001110100010 : VALUE=19'b0000000_101010111001;
      15'b010_001110100011 : VALUE=19'b0000000_101010111001;
      15'b010_001110100100 : VALUE=19'b0000000_101010111000;
      15'b010_001110100101 : VALUE=19'b0000000_101010111000;
      15'b010_001110100110 : VALUE=19'b0000000_101010111000;
      15'b010_001110100111 : VALUE=19'b0000000_101010111000;
      15'b010_001110101000 : VALUE=19'b0000000_101010111000;
      15'b010_001110101001 : VALUE=19'b0000000_101010111000;
      15'b010_001110101010 : VALUE=19'b0000000_101010110111;
      15'b010_001110101011 : VALUE=19'b0000000_101010110111;
      15'b010_001110101100 : VALUE=19'b0000000_101010110111;
      15'b010_001110101101 : VALUE=19'b0000000_101010110111;
      15'b010_001110101110 : VALUE=19'b0000000_101010110111;
      15'b010_001110101111 : VALUE=19'b0000000_101010110111;
      15'b010_001110110000 : VALUE=19'b0000000_101010110111;
      15'b010_001110110001 : VALUE=19'b0000000_101010110110;
      15'b010_001110110010 : VALUE=19'b0000000_101010110110;
      15'b010_001110110011 : VALUE=19'b0000000_101010110110;
      15'b010_001110110100 : VALUE=19'b0000000_101010110110;
      15'b010_001110110101 : VALUE=19'b0000000_101010110110;
      15'b010_001110110110 : VALUE=19'b0000000_101010110110;
      15'b010_001110110111 : VALUE=19'b0000000_101010110110;
      15'b010_001110111000 : VALUE=19'b0000000_101010110101;
      15'b010_001110111001 : VALUE=19'b0000000_101010110101;
      15'b010_001110111010 : VALUE=19'b0000000_101010110101;
      15'b010_001110111011 : VALUE=19'b0000000_101010110101;
      15'b010_001110111100 : VALUE=19'b0000000_101010110101;
      15'b010_001110111101 : VALUE=19'b0000000_101010110101;
      15'b010_001110111110 : VALUE=19'b0000000_101010110100;
      15'b010_001110111111 : VALUE=19'b0000000_101010110100;
      15'b010_001111000000 : VALUE=19'b0000000_101010110100;
      15'b010_001111000001 : VALUE=19'b0000000_101010110100;
      15'b010_001111000010 : VALUE=19'b0000000_101010110100;
      15'b010_001111000011 : VALUE=19'b0000000_101010110100;
      15'b010_001111000100 : VALUE=19'b0000000_101010110100;
      15'b010_001111000101 : VALUE=19'b0000000_101010110011;
      15'b010_001111000110 : VALUE=19'b0000000_101010110011;
      15'b010_001111000111 : VALUE=19'b0000000_101010110011;
      15'b010_001111001000 : VALUE=19'b0000000_101010110011;
      15'b010_001111001001 : VALUE=19'b0000000_101010110011;
      15'b010_001111001010 : VALUE=19'b0000000_101010110011;
      15'b010_001111001011 : VALUE=19'b0000000_101010110011;
      15'b010_001111001100 : VALUE=19'b0000000_101010110010;
      15'b010_001111001101 : VALUE=19'b0000000_101010110010;
      15'b010_001111001110 : VALUE=19'b0000000_101010110010;
      15'b010_001111001111 : VALUE=19'b0000000_101010110010;
      15'b010_001111010000 : VALUE=19'b0000000_101010110010;
      15'b010_001111010001 : VALUE=19'b0000000_101010110010;
      15'b010_001111010010 : VALUE=19'b0000000_101010110010;
      15'b010_001111010011 : VALUE=19'b0000000_101010110001;
      15'b010_001111010100 : VALUE=19'b0000000_101010110001;
      15'b010_001111010101 : VALUE=19'b0000000_101010110001;
      15'b010_001111010110 : VALUE=19'b0000000_101010110001;
      15'b010_001111010111 : VALUE=19'b0000000_101010110001;
      15'b010_001111011000 : VALUE=19'b0000000_101010110001;
      15'b010_001111011001 : VALUE=19'b0000000_101010110000;
      15'b010_001111011010 : VALUE=19'b0000000_101010110000;
      15'b010_001111011011 : VALUE=19'b0000000_101010110000;
      15'b010_001111011100 : VALUE=19'b0000000_101010110000;
      15'b010_001111011101 : VALUE=19'b0000000_101010110000;
      15'b010_001111011110 : VALUE=19'b0000000_101010110000;
      15'b010_001111011111 : VALUE=19'b0000000_101010110000;
      15'b010_001111100000 : VALUE=19'b0000000_101010101111;
      15'b010_001111100001 : VALUE=19'b0000000_101010101111;
      15'b010_001111100010 : VALUE=19'b0000000_101010101111;
      15'b010_001111100011 : VALUE=19'b0000000_101010101111;
      15'b010_001111100100 : VALUE=19'b0000000_101010101111;
      15'b010_001111100101 : VALUE=19'b0000000_101010101111;
      15'b010_001111100110 : VALUE=19'b0000000_101010101111;
      15'b010_001111100111 : VALUE=19'b0000000_101010101110;
      15'b010_001111101000 : VALUE=19'b0000000_101010101110;
      15'b010_001111101001 : VALUE=19'b0000000_101010101110;
      15'b010_001111101010 : VALUE=19'b0000000_101010101110;
      15'b010_001111101011 : VALUE=19'b0000000_101010101110;
      15'b010_001111101100 : VALUE=19'b0000000_101010101110;
      15'b010_001111101101 : VALUE=19'b0000000_101010101101;
      15'b010_001111101110 : VALUE=19'b0000000_101010101101;
      15'b010_001111101111 : VALUE=19'b0000000_101010101101;
      15'b010_001111110000 : VALUE=19'b0000000_101010101101;
      15'b010_001111110001 : VALUE=19'b0000000_101010101101;
      15'b010_001111110010 : VALUE=19'b0000000_101010101101;
      15'b010_001111110011 : VALUE=19'b0000000_101010101101;
      15'b010_001111110100 : VALUE=19'b0000000_101010101100;
      15'b010_001111110101 : VALUE=19'b0000000_101010101100;
      15'b010_001111110110 : VALUE=19'b0000000_101010101100;
      15'b010_001111110111 : VALUE=19'b0000000_101010101100;
      15'b010_001111111000 : VALUE=19'b0000000_101010101100;
      15'b010_001111111001 : VALUE=19'b0000000_101010101100;
      15'b010_001111111010 : VALUE=19'b0000000_101010101100;
      15'b010_001111111011 : VALUE=19'b0000000_101010101011;
      15'b010_001111111100 : VALUE=19'b0000000_101010101011;
      15'b010_001111111101 : VALUE=19'b0000000_101010101011;
      15'b010_001111111110 : VALUE=19'b0000000_101010101011;
      15'b010_001111111111 : VALUE=19'b0000000_101010101011;
      15'b010_010000000000 : VALUE=19'b0000000_101010101011;
      15'b010_010000000001 : VALUE=19'b0000000_101010101011;
      15'b010_010000000010 : VALUE=19'b0000000_101010101010;
      15'b010_010000000011 : VALUE=19'b0000000_101010101010;
      15'b010_010000000100 : VALUE=19'b0000000_101010101010;
      15'b010_010000000101 : VALUE=19'b0000000_101010101010;
      15'b010_010000000110 : VALUE=19'b0000000_101010101010;
      15'b010_010000000111 : VALUE=19'b0000000_101010101010;
      15'b010_010000001000 : VALUE=19'b0000000_101010101001;
      15'b010_010000001001 : VALUE=19'b0000000_101010101001;
      15'b010_010000001010 : VALUE=19'b0000000_101010101001;
      15'b010_010000001011 : VALUE=19'b0000000_101010101001;
      15'b010_010000001100 : VALUE=19'b0000000_101010101001;
      15'b010_010000001101 : VALUE=19'b0000000_101010101001;
      15'b010_010000001110 : VALUE=19'b0000000_101010101001;
      15'b010_010000001111 : VALUE=19'b0000000_101010101000;
      15'b010_010000010000 : VALUE=19'b0000000_101010101000;
      15'b010_010000010001 : VALUE=19'b0000000_101010101000;
      15'b010_010000010010 : VALUE=19'b0000000_101010101000;
      15'b010_010000010011 : VALUE=19'b0000000_101010101000;
      15'b010_010000010100 : VALUE=19'b0000000_101010101000;
      15'b010_010000010101 : VALUE=19'b0000000_101010101000;
      15'b010_010000010110 : VALUE=19'b0000000_101010100111;
      15'b010_010000010111 : VALUE=19'b0000000_101010100111;
      15'b010_010000011000 : VALUE=19'b0000000_101010100111;
      15'b010_010000011001 : VALUE=19'b0000000_101010100111;
      15'b010_010000011010 : VALUE=19'b0000000_101010100111;
      15'b010_010000011011 : VALUE=19'b0000000_101010100111;
      15'b010_010000011100 : VALUE=19'b0000000_101010100111;
      15'b010_010000011101 : VALUE=19'b0000000_101010100110;
      15'b010_010000011110 : VALUE=19'b0000000_101010100110;
      15'b010_010000011111 : VALUE=19'b0000000_101010100110;
      15'b010_010000100000 : VALUE=19'b0000000_101010100110;
      15'b010_010000100001 : VALUE=19'b0000000_101010100110;
      15'b010_010000100010 : VALUE=19'b0000000_101010100110;
      15'b010_010000100011 : VALUE=19'b0000000_101010100101;
      15'b010_010000100100 : VALUE=19'b0000000_101010100101;
      15'b010_010000100101 : VALUE=19'b0000000_101010100101;
      15'b010_010000100110 : VALUE=19'b0000000_101010100101;
      15'b010_010000100111 : VALUE=19'b0000000_101010100101;
      15'b010_010000101000 : VALUE=19'b0000000_101010100101;
      15'b010_010000101001 : VALUE=19'b0000000_101010100101;
      15'b010_010000101010 : VALUE=19'b0000000_101010100100;
      15'b010_010000101011 : VALUE=19'b0000000_101010100100;
      15'b010_010000101100 : VALUE=19'b0000000_101010100100;
      15'b010_010000101101 : VALUE=19'b0000000_101010100100;
      15'b010_010000101110 : VALUE=19'b0000000_101010100100;
      15'b010_010000101111 : VALUE=19'b0000000_101010100100;
      15'b010_010000110000 : VALUE=19'b0000000_101010100100;
      15'b010_010000110001 : VALUE=19'b0000000_101010100011;
      15'b010_010000110010 : VALUE=19'b0000000_101010100011;
      15'b010_010000110011 : VALUE=19'b0000000_101010100011;
      15'b010_010000110100 : VALUE=19'b0000000_101010100011;
      15'b010_010000110101 : VALUE=19'b0000000_101010100011;
      15'b010_010000110110 : VALUE=19'b0000000_101010100011;
      15'b010_010000110111 : VALUE=19'b0000000_101010100011;
      15'b010_010000111000 : VALUE=19'b0000000_101010100010;
      15'b010_010000111001 : VALUE=19'b0000000_101010100010;
      15'b010_010000111010 : VALUE=19'b0000000_101010100010;
      15'b010_010000111011 : VALUE=19'b0000000_101010100010;
      15'b010_010000111100 : VALUE=19'b0000000_101010100010;
      15'b010_010000111101 : VALUE=19'b0000000_101010100010;
      15'b010_010000111110 : VALUE=19'b0000000_101010100010;
      15'b010_010000111111 : VALUE=19'b0000000_101010100001;
      15'b010_010001000000 : VALUE=19'b0000000_101010100001;
      15'b010_010001000001 : VALUE=19'b0000000_101010100001;
      15'b010_010001000010 : VALUE=19'b0000000_101010100001;
      15'b010_010001000011 : VALUE=19'b0000000_101010100001;
      15'b010_010001000100 : VALUE=19'b0000000_101010100001;
      15'b010_010001000101 : VALUE=19'b0000000_101010100001;
      15'b010_010001000110 : VALUE=19'b0000000_101010100000;
      15'b010_010001000111 : VALUE=19'b0000000_101010100000;
      15'b010_010001001000 : VALUE=19'b0000000_101010100000;
      15'b010_010001001001 : VALUE=19'b0000000_101010100000;
      15'b010_010001001010 : VALUE=19'b0000000_101010100000;
      15'b010_010001001011 : VALUE=19'b0000000_101010100000;
      15'b010_010001001100 : VALUE=19'b0000000_101010011111;
      15'b010_010001001101 : VALUE=19'b0000000_101010011111;
      15'b010_010001001110 : VALUE=19'b0000000_101010011111;
      15'b010_010001001111 : VALUE=19'b0000000_101010011111;
      15'b010_010001010000 : VALUE=19'b0000000_101010011111;
      15'b010_010001010001 : VALUE=19'b0000000_101010011111;
      15'b010_010001010010 : VALUE=19'b0000000_101010011111;
      15'b010_010001010011 : VALUE=19'b0000000_101010011110;
      15'b010_010001010100 : VALUE=19'b0000000_101010011110;
      15'b010_010001010101 : VALUE=19'b0000000_101010011110;
      15'b010_010001010110 : VALUE=19'b0000000_101010011110;
      15'b010_010001010111 : VALUE=19'b0000000_101010011110;
      15'b010_010001011000 : VALUE=19'b0000000_101010011110;
      15'b010_010001011001 : VALUE=19'b0000000_101010011110;
      15'b010_010001011010 : VALUE=19'b0000000_101010011101;
      15'b010_010001011011 : VALUE=19'b0000000_101010011101;
      15'b010_010001011100 : VALUE=19'b0000000_101010011101;
      15'b010_010001011101 : VALUE=19'b0000000_101010011101;
      15'b010_010001011110 : VALUE=19'b0000000_101010011101;
      15'b010_010001011111 : VALUE=19'b0000000_101010011101;
      15'b010_010001100000 : VALUE=19'b0000000_101010011101;
      15'b010_010001100001 : VALUE=19'b0000000_101010011100;
      15'b010_010001100010 : VALUE=19'b0000000_101010011100;
      15'b010_010001100011 : VALUE=19'b0000000_101010011100;
      15'b010_010001100100 : VALUE=19'b0000000_101010011100;
      15'b010_010001100101 : VALUE=19'b0000000_101010011100;
      15'b010_010001100110 : VALUE=19'b0000000_101010011100;
      15'b010_010001100111 : VALUE=19'b0000000_101010011100;
      15'b010_010001101000 : VALUE=19'b0000000_101010011011;
      15'b010_010001101001 : VALUE=19'b0000000_101010011011;
      15'b010_010001101010 : VALUE=19'b0000000_101010011011;
      15'b010_010001101011 : VALUE=19'b0000000_101010011011;
      15'b010_010001101100 : VALUE=19'b0000000_101010011011;
      15'b010_010001101101 : VALUE=19'b0000000_101010011011;
      15'b010_010001101110 : VALUE=19'b0000000_101010011011;
      15'b010_010001101111 : VALUE=19'b0000000_101010011010;
      15'b010_010001110000 : VALUE=19'b0000000_101010011010;
      15'b010_010001110001 : VALUE=19'b0000000_101010011010;
      15'b010_010001110010 : VALUE=19'b0000000_101010011010;
      15'b010_010001110011 : VALUE=19'b0000000_101010011010;
      15'b010_010001110100 : VALUE=19'b0000000_101010011010;
      15'b010_010001110101 : VALUE=19'b0000000_101010011001;
      15'b010_010001110110 : VALUE=19'b0000000_101010011001;
      15'b010_010001110111 : VALUE=19'b0000000_101010011001;
      15'b010_010001111000 : VALUE=19'b0000000_101010011001;
      15'b010_010001111001 : VALUE=19'b0000000_101010011001;
      15'b010_010001111010 : VALUE=19'b0000000_101010011001;
      15'b010_010001111011 : VALUE=19'b0000000_101010011001;
      15'b010_010001111100 : VALUE=19'b0000000_101010011000;
      15'b010_010001111101 : VALUE=19'b0000000_101010011000;
      15'b010_010001111110 : VALUE=19'b0000000_101010011000;
      15'b010_010001111111 : VALUE=19'b0000000_101010011000;
      15'b010_010010000000 : VALUE=19'b0000000_101010011000;
      15'b010_010010000001 : VALUE=19'b0000000_101010011000;
      15'b010_010010000010 : VALUE=19'b0000000_101010011000;
      15'b010_010010000011 : VALUE=19'b0000000_101010010111;
      15'b010_010010000100 : VALUE=19'b0000000_101010010111;
      15'b010_010010000101 : VALUE=19'b0000000_101010010111;
      15'b010_010010000110 : VALUE=19'b0000000_101010010111;
      15'b010_010010000111 : VALUE=19'b0000000_101010010111;
      15'b010_010010001000 : VALUE=19'b0000000_101010010111;
      15'b010_010010001001 : VALUE=19'b0000000_101010010111;
      15'b010_010010001010 : VALUE=19'b0000000_101010010110;
      15'b010_010010001011 : VALUE=19'b0000000_101010010110;
      15'b010_010010001100 : VALUE=19'b0000000_101010010110;
      15'b010_010010001101 : VALUE=19'b0000000_101010010110;
      15'b010_010010001110 : VALUE=19'b0000000_101010010110;
      15'b010_010010001111 : VALUE=19'b0000000_101010010110;
      15'b010_010010010000 : VALUE=19'b0000000_101010010110;
      15'b010_010010010001 : VALUE=19'b0000000_101010010101;
      15'b010_010010010010 : VALUE=19'b0000000_101010010101;
      15'b010_010010010011 : VALUE=19'b0000000_101010010101;
      15'b010_010010010100 : VALUE=19'b0000000_101010010101;
      15'b010_010010010101 : VALUE=19'b0000000_101010010101;
      15'b010_010010010110 : VALUE=19'b0000000_101010010101;
      15'b010_010010010111 : VALUE=19'b0000000_101010010101;
      15'b010_010010011000 : VALUE=19'b0000000_101010010100;
      15'b010_010010011001 : VALUE=19'b0000000_101010010100;
      15'b010_010010011010 : VALUE=19'b0000000_101010010100;
      15'b010_010010011011 : VALUE=19'b0000000_101010010100;
      15'b010_010010011100 : VALUE=19'b0000000_101010010100;
      15'b010_010010011101 : VALUE=19'b0000000_101010010100;
      15'b010_010010011110 : VALUE=19'b0000000_101010010100;
      15'b010_010010011111 : VALUE=19'b0000000_101010010011;
      15'b010_010010100000 : VALUE=19'b0000000_101010010011;
      15'b010_010010100001 : VALUE=19'b0000000_101010010011;
      15'b010_010010100010 : VALUE=19'b0000000_101010010011;
      15'b010_010010100011 : VALUE=19'b0000000_101010010011;
      15'b010_010010100100 : VALUE=19'b0000000_101010010011;
      15'b010_010010100101 : VALUE=19'b0000000_101010010011;
      15'b010_010010100110 : VALUE=19'b0000000_101010010010;
      15'b010_010010100111 : VALUE=19'b0000000_101010010010;
      15'b010_010010101000 : VALUE=19'b0000000_101010010010;
      15'b010_010010101001 : VALUE=19'b0000000_101010010010;
      15'b010_010010101010 : VALUE=19'b0000000_101010010010;
      15'b010_010010101011 : VALUE=19'b0000000_101010010010;
      15'b010_010010101100 : VALUE=19'b0000000_101010010010;
      15'b010_010010101101 : VALUE=19'b0000000_101010010001;
      15'b010_010010101110 : VALUE=19'b0000000_101010010001;
      15'b010_010010101111 : VALUE=19'b0000000_101010010001;
      15'b010_010010110000 : VALUE=19'b0000000_101010010001;
      15'b010_010010110001 : VALUE=19'b0000000_101010010001;
      15'b010_010010110010 : VALUE=19'b0000000_101010010001;
      15'b010_010010110011 : VALUE=19'b0000000_101010010001;
      15'b010_010010110100 : VALUE=19'b0000000_101010010000;
      15'b010_010010110101 : VALUE=19'b0000000_101010010000;
      15'b010_010010110110 : VALUE=19'b0000000_101010010000;
      15'b010_010010110111 : VALUE=19'b0000000_101010010000;
      15'b010_010010111000 : VALUE=19'b0000000_101010010000;
      15'b010_010010111001 : VALUE=19'b0000000_101010010000;
      15'b010_010010111010 : VALUE=19'b0000000_101010010000;
      15'b010_010010111011 : VALUE=19'b0000000_101010001111;
      15'b010_010010111100 : VALUE=19'b0000000_101010001111;
      15'b010_010010111101 : VALUE=19'b0000000_101010001111;
      15'b010_010010111110 : VALUE=19'b0000000_101010001111;
      15'b010_010010111111 : VALUE=19'b0000000_101010001111;
      15'b010_010011000000 : VALUE=19'b0000000_101010001111;
      15'b010_010011000001 : VALUE=19'b0000000_101010001111;
      15'b010_010011000010 : VALUE=19'b0000000_101010001110;
      15'b010_010011000011 : VALUE=19'b0000000_101010001110;
      15'b010_010011000100 : VALUE=19'b0000000_101010001110;
      15'b010_010011000101 : VALUE=19'b0000000_101010001110;
      15'b010_010011000110 : VALUE=19'b0000000_101010001110;
      15'b010_010011000111 : VALUE=19'b0000000_101010001110;
      15'b010_010011001000 : VALUE=19'b0000000_101010001110;
      15'b010_010011001001 : VALUE=19'b0000000_101010001101;
      15'b010_010011001010 : VALUE=19'b0000000_101010001101;
      15'b010_010011001011 : VALUE=19'b0000000_101010001101;
      15'b010_010011001100 : VALUE=19'b0000000_101010001101;
      15'b010_010011001101 : VALUE=19'b0000000_101010001101;
      15'b010_010011001110 : VALUE=19'b0000000_101010001101;
      15'b010_010011001111 : VALUE=19'b0000000_101010001101;
      15'b010_010011010000 : VALUE=19'b0000000_101010001100;
      15'b010_010011010001 : VALUE=19'b0000000_101010001100;
      15'b010_010011010010 : VALUE=19'b0000000_101010001100;
      15'b010_010011010011 : VALUE=19'b0000000_101010001100;
      15'b010_010011010100 : VALUE=19'b0000000_101010001100;
      15'b010_010011010101 : VALUE=19'b0000000_101010001100;
      15'b010_010011010110 : VALUE=19'b0000000_101010001100;
      15'b010_010011010111 : VALUE=19'b0000000_101010001011;
      15'b010_010011011000 : VALUE=19'b0000000_101010001011;
      15'b010_010011011001 : VALUE=19'b0000000_101010001011;
      15'b010_010011011010 : VALUE=19'b0000000_101010001011;
      15'b010_010011011011 : VALUE=19'b0000000_101010001011;
      15'b010_010011011100 : VALUE=19'b0000000_101010001011;
      15'b010_010011011101 : VALUE=19'b0000000_101010001011;
      15'b010_010011011110 : VALUE=19'b0000000_101010001010;
      15'b010_010011011111 : VALUE=19'b0000000_101010001010;
      15'b010_010011100000 : VALUE=19'b0000000_101010001010;
      15'b010_010011100001 : VALUE=19'b0000000_101010001010;
      15'b010_010011100010 : VALUE=19'b0000000_101010001010;
      15'b010_010011100011 : VALUE=19'b0000000_101010001010;
      15'b010_010011100100 : VALUE=19'b0000000_101010001010;
      15'b010_010011100101 : VALUE=19'b0000000_101010001001;
      15'b010_010011100110 : VALUE=19'b0000000_101010001001;
      15'b010_010011100111 : VALUE=19'b0000000_101010001001;
      15'b010_010011101000 : VALUE=19'b0000000_101010001001;
      15'b010_010011101001 : VALUE=19'b0000000_101010001001;
      15'b010_010011101010 : VALUE=19'b0000000_101010001001;
      15'b010_010011101011 : VALUE=19'b0000000_101010001001;
      15'b010_010011101100 : VALUE=19'b0000000_101010001000;
      15'b010_010011101101 : VALUE=19'b0000000_101010001000;
      15'b010_010011101110 : VALUE=19'b0000000_101010001000;
      15'b010_010011101111 : VALUE=19'b0000000_101010001000;
      15'b010_010011110000 : VALUE=19'b0000000_101010001000;
      15'b010_010011110001 : VALUE=19'b0000000_101010001000;
      15'b010_010011110010 : VALUE=19'b0000000_101010001000;
      15'b010_010011110011 : VALUE=19'b0000000_101010000111;
      15'b010_010011110100 : VALUE=19'b0000000_101010000111;
      15'b010_010011110101 : VALUE=19'b0000000_101010000111;
      15'b010_010011110110 : VALUE=19'b0000000_101010000111;
      15'b010_010011110111 : VALUE=19'b0000000_101010000111;
      15'b010_010011111000 : VALUE=19'b0000000_101010000111;
      15'b010_010011111001 : VALUE=19'b0000000_101010000111;
      15'b010_010011111010 : VALUE=19'b0000000_101010000110;
      15'b010_010011111011 : VALUE=19'b0000000_101010000110;
      15'b010_010011111100 : VALUE=19'b0000000_101010000110;
      15'b010_010011111101 : VALUE=19'b0000000_101010000110;
      15'b010_010011111110 : VALUE=19'b0000000_101010000110;
      15'b010_010011111111 : VALUE=19'b0000000_101010000110;
      15'b010_010100000000 : VALUE=19'b0000000_101010000110;
      15'b010_010100000001 : VALUE=19'b0000000_101010000101;
      15'b010_010100000010 : VALUE=19'b0000000_101010000101;
      15'b010_010100000011 : VALUE=19'b0000000_101010000101;
      15'b010_010100000100 : VALUE=19'b0000000_101010000101;
      15'b010_010100000101 : VALUE=19'b0000000_101010000101;
      15'b010_010100000110 : VALUE=19'b0000000_101010000101;
      15'b010_010100000111 : VALUE=19'b0000000_101010000101;
      15'b010_010100001000 : VALUE=19'b0000000_101010000100;
      15'b010_010100001001 : VALUE=19'b0000000_101010000100;
      15'b010_010100001010 : VALUE=19'b0000000_101010000100;
      15'b010_010100001011 : VALUE=19'b0000000_101010000100;
      15'b010_010100001100 : VALUE=19'b0000000_101010000100;
      15'b010_010100001101 : VALUE=19'b0000000_101010000100;
      15'b010_010100001110 : VALUE=19'b0000000_101010000100;
      15'b010_010100001111 : VALUE=19'b0000000_101010000011;
      15'b010_010100010000 : VALUE=19'b0000000_101010000011;
      15'b010_010100010001 : VALUE=19'b0000000_101010000011;
      15'b010_010100010010 : VALUE=19'b0000000_101010000011;
      15'b010_010100010011 : VALUE=19'b0000000_101010000011;
      15'b010_010100010100 : VALUE=19'b0000000_101010000011;
      15'b010_010100010101 : VALUE=19'b0000000_101010000011;
      15'b010_010100010110 : VALUE=19'b0000000_101010000010;
      15'b010_010100010111 : VALUE=19'b0000000_101010000010;
      15'b010_010100011000 : VALUE=19'b0000000_101010000010;
      15'b010_010100011001 : VALUE=19'b0000000_101010000010;
      15'b010_010100011010 : VALUE=19'b0000000_101010000010;
      15'b010_010100011011 : VALUE=19'b0000000_101010000010;
      15'b010_010100011100 : VALUE=19'b0000000_101010000010;
      15'b010_010100011101 : VALUE=19'b0000000_101010000001;
      15'b010_010100011110 : VALUE=19'b0000000_101010000001;
      15'b010_010100011111 : VALUE=19'b0000000_101010000001;
      15'b010_010100100000 : VALUE=19'b0000000_101010000001;
      15'b010_010100100001 : VALUE=19'b0000000_101010000001;
      15'b010_010100100010 : VALUE=19'b0000000_101010000001;
      15'b010_010100100011 : VALUE=19'b0000000_101010000001;
      15'b010_010100100100 : VALUE=19'b0000000_101010000000;
      15'b010_010100100101 : VALUE=19'b0000000_101010000000;
      15'b010_010100100110 : VALUE=19'b0000000_101010000000;
      15'b010_010100100111 : VALUE=19'b0000000_101010000000;
      15'b010_010100101000 : VALUE=19'b0000000_101010000000;
      15'b010_010100101001 : VALUE=19'b0000000_101010000000;
      15'b010_010100101010 : VALUE=19'b0000000_101010000000;
      15'b010_010100101011 : VALUE=19'b0000000_101001111111;
      15'b010_010100101100 : VALUE=19'b0000000_101001111111;
      15'b010_010100101101 : VALUE=19'b0000000_101001111111;
      15'b010_010100101110 : VALUE=19'b0000000_101001111111;
      15'b010_010100101111 : VALUE=19'b0000000_101001111111;
      15'b010_010100110000 : VALUE=19'b0000000_101001111111;
      15'b010_010100110001 : VALUE=19'b0000000_101001111111;
      15'b010_010100110010 : VALUE=19'b0000000_101001111110;
      15'b010_010100110011 : VALUE=19'b0000000_101001111110;
      15'b010_010100110100 : VALUE=19'b0000000_101001111110;
      15'b010_010100110101 : VALUE=19'b0000000_101001111110;
      15'b010_010100110110 : VALUE=19'b0000000_101001111110;
      15'b010_010100110111 : VALUE=19'b0000000_101001111110;
      15'b010_010100111000 : VALUE=19'b0000000_101001111110;
      15'b010_010100111001 : VALUE=19'b0000000_101001111101;
      15'b010_010100111010 : VALUE=19'b0000000_101001111101;
      15'b010_010100111011 : VALUE=19'b0000000_101001111101;
      15'b010_010100111100 : VALUE=19'b0000000_101001111101;
      15'b010_010100111101 : VALUE=19'b0000000_101001111101;
      15'b010_010100111110 : VALUE=19'b0000000_101001111101;
      15'b010_010100111111 : VALUE=19'b0000000_101001111101;
      15'b010_010101000000 : VALUE=19'b0000000_101001111100;
      15'b010_010101000001 : VALUE=19'b0000000_101001111100;
      15'b010_010101000010 : VALUE=19'b0000000_101001111100;
      15'b010_010101000011 : VALUE=19'b0000000_101001111100;
      15'b010_010101000100 : VALUE=19'b0000000_101001111100;
      15'b010_010101000101 : VALUE=19'b0000000_101001111100;
      15'b010_010101000110 : VALUE=19'b0000000_101001111100;
      15'b010_010101000111 : VALUE=19'b0000000_101001111011;
      15'b010_010101001000 : VALUE=19'b0000000_101001111011;
      15'b010_010101001001 : VALUE=19'b0000000_101001111011;
      15'b010_010101001010 : VALUE=19'b0000000_101001111011;
      15'b010_010101001011 : VALUE=19'b0000000_101001111011;
      15'b010_010101001100 : VALUE=19'b0000000_101001111011;
      15'b010_010101001101 : VALUE=19'b0000000_101001111011;
      15'b010_010101001110 : VALUE=19'b0000000_101001111010;
      15'b010_010101001111 : VALUE=19'b0000000_101001111010;
      15'b010_010101010000 : VALUE=19'b0000000_101001111010;
      15'b010_010101010001 : VALUE=19'b0000000_101001111010;
      15'b010_010101010010 : VALUE=19'b0000000_101001111010;
      15'b010_010101010011 : VALUE=19'b0000000_101001111010;
      15'b010_010101010100 : VALUE=19'b0000000_101001111010;
      15'b010_010101010101 : VALUE=19'b0000000_101001111010;
      15'b010_010101010110 : VALUE=19'b0000000_101001111001;
      15'b010_010101010111 : VALUE=19'b0000000_101001111001;
      15'b010_010101011000 : VALUE=19'b0000000_101001111001;
      15'b010_010101011001 : VALUE=19'b0000000_101001111001;
      15'b010_010101011010 : VALUE=19'b0000000_101001111001;
      15'b010_010101011011 : VALUE=19'b0000000_101001111001;
      15'b010_010101011100 : VALUE=19'b0000000_101001111001;
      15'b010_010101011101 : VALUE=19'b0000000_101001111000;
      15'b010_010101011110 : VALUE=19'b0000000_101001111000;
      15'b010_010101011111 : VALUE=19'b0000000_101001111000;
      15'b010_010101100000 : VALUE=19'b0000000_101001111000;
      15'b010_010101100001 : VALUE=19'b0000000_101001111000;
      15'b010_010101100010 : VALUE=19'b0000000_101001111000;
      15'b010_010101100011 : VALUE=19'b0000000_101001111000;
      15'b010_010101100100 : VALUE=19'b0000000_101001110111;
      15'b010_010101100101 : VALUE=19'b0000000_101001110111;
      15'b010_010101100110 : VALUE=19'b0000000_101001110111;
      15'b010_010101100111 : VALUE=19'b0000000_101001110111;
      15'b010_010101101000 : VALUE=19'b0000000_101001110111;
      15'b010_010101101001 : VALUE=19'b0000000_101001110111;
      15'b010_010101101010 : VALUE=19'b0000000_101001110111;
      15'b010_010101101011 : VALUE=19'b0000000_101001110110;
      15'b010_010101101100 : VALUE=19'b0000000_101001110110;
      15'b010_010101101101 : VALUE=19'b0000000_101001110110;
      15'b010_010101101110 : VALUE=19'b0000000_101001110110;
      15'b010_010101101111 : VALUE=19'b0000000_101001110110;
      15'b010_010101110000 : VALUE=19'b0000000_101001110110;
      15'b010_010101110001 : VALUE=19'b0000000_101001110110;
      15'b010_010101110010 : VALUE=19'b0000000_101001110101;
      15'b010_010101110011 : VALUE=19'b0000000_101001110101;
      15'b010_010101110100 : VALUE=19'b0000000_101001110101;
      15'b010_010101110101 : VALUE=19'b0000000_101001110101;
      15'b010_010101110110 : VALUE=19'b0000000_101001110101;
      15'b010_010101110111 : VALUE=19'b0000000_101001110101;
      15'b010_010101111000 : VALUE=19'b0000000_101001110101;
      15'b010_010101111001 : VALUE=19'b0000000_101001110100;
      15'b010_010101111010 : VALUE=19'b0000000_101001110100;
      15'b010_010101111011 : VALUE=19'b0000000_101001110100;
      15'b010_010101111100 : VALUE=19'b0000000_101001110100;
      15'b010_010101111101 : VALUE=19'b0000000_101001110100;
      15'b010_010101111110 : VALUE=19'b0000000_101001110100;
      15'b010_010101111111 : VALUE=19'b0000000_101001110100;
      15'b010_010110000000 : VALUE=19'b0000000_101001110011;
      15'b010_010110000001 : VALUE=19'b0000000_101001110011;
      15'b010_010110000010 : VALUE=19'b0000000_101001110011;
      15'b010_010110000011 : VALUE=19'b0000000_101001110011;
      15'b010_010110000100 : VALUE=19'b0000000_101001110011;
      15'b010_010110000101 : VALUE=19'b0000000_101001110011;
      15'b010_010110000110 : VALUE=19'b0000000_101001110011;
      15'b010_010110000111 : VALUE=19'b0000000_101001110011;
      15'b010_010110001000 : VALUE=19'b0000000_101001110010;
      15'b010_010110001001 : VALUE=19'b0000000_101001110010;
      15'b010_010110001010 : VALUE=19'b0000000_101001110010;
      15'b010_010110001011 : VALUE=19'b0000000_101001110010;
      15'b010_010110001100 : VALUE=19'b0000000_101001110010;
      15'b010_010110001101 : VALUE=19'b0000000_101001110010;
      15'b010_010110001110 : VALUE=19'b0000000_101001110010;
      15'b010_010110001111 : VALUE=19'b0000000_101001110001;
      15'b010_010110010000 : VALUE=19'b0000000_101001110001;
      15'b010_010110010001 : VALUE=19'b0000000_101001110001;
      15'b010_010110010010 : VALUE=19'b0000000_101001110001;
      15'b010_010110010011 : VALUE=19'b0000000_101001110001;
      15'b010_010110010100 : VALUE=19'b0000000_101001110001;
      15'b010_010110010101 : VALUE=19'b0000000_101001110001;
      15'b010_010110010110 : VALUE=19'b0000000_101001110000;
      15'b010_010110010111 : VALUE=19'b0000000_101001110000;
      15'b010_010110011000 : VALUE=19'b0000000_101001110000;
      15'b010_010110011001 : VALUE=19'b0000000_101001110000;
      15'b010_010110011010 : VALUE=19'b0000000_101001110000;
      15'b010_010110011011 : VALUE=19'b0000000_101001110000;
      15'b010_010110011100 : VALUE=19'b0000000_101001110000;
      15'b010_010110011101 : VALUE=19'b0000000_101001101111;
      15'b010_010110011110 : VALUE=19'b0000000_101001101111;
      15'b010_010110011111 : VALUE=19'b0000000_101001101111;
      15'b010_010110100000 : VALUE=19'b0000000_101001101111;
      15'b010_010110100001 : VALUE=19'b0000000_101001101111;
      15'b010_010110100010 : VALUE=19'b0000000_101001101111;
      15'b010_010110100011 : VALUE=19'b0000000_101001101111;
      15'b010_010110100100 : VALUE=19'b0000000_101001101110;
      15'b010_010110100101 : VALUE=19'b0000000_101001101110;
      15'b010_010110100110 : VALUE=19'b0000000_101001101110;
      15'b010_010110100111 : VALUE=19'b0000000_101001101110;
      15'b010_010110101000 : VALUE=19'b0000000_101001101110;
      15'b010_010110101001 : VALUE=19'b0000000_101001101110;
      15'b010_010110101010 : VALUE=19'b0000000_101001101110;
      15'b010_010110101011 : VALUE=19'b0000000_101001101110;
      15'b010_010110101100 : VALUE=19'b0000000_101001101101;
      15'b010_010110101101 : VALUE=19'b0000000_101001101101;
      15'b010_010110101110 : VALUE=19'b0000000_101001101101;
      15'b010_010110101111 : VALUE=19'b0000000_101001101101;
      15'b010_010110110000 : VALUE=19'b0000000_101001101101;
      15'b010_010110110001 : VALUE=19'b0000000_101001101101;
      15'b010_010110110010 : VALUE=19'b0000000_101001101101;
      15'b010_010110110011 : VALUE=19'b0000000_101001101100;
      15'b010_010110110100 : VALUE=19'b0000000_101001101100;
      15'b010_010110110101 : VALUE=19'b0000000_101001101100;
      15'b010_010110110110 : VALUE=19'b0000000_101001101100;
      15'b010_010110110111 : VALUE=19'b0000000_101001101100;
      15'b010_010110111000 : VALUE=19'b0000000_101001101100;
      15'b010_010110111001 : VALUE=19'b0000000_101001101100;
      15'b010_010110111010 : VALUE=19'b0000000_101001101011;
      15'b010_010110111011 : VALUE=19'b0000000_101001101011;
      15'b010_010110111100 : VALUE=19'b0000000_101001101011;
      15'b010_010110111101 : VALUE=19'b0000000_101001101011;
      15'b010_010110111110 : VALUE=19'b0000000_101001101011;
      15'b010_010110111111 : VALUE=19'b0000000_101001101011;
      15'b010_010111000000 : VALUE=19'b0000000_101001101011;
      15'b010_010111000001 : VALUE=19'b0000000_101001101010;
      15'b010_010111000010 : VALUE=19'b0000000_101001101010;
      15'b010_010111000011 : VALUE=19'b0000000_101001101010;
      15'b010_010111000100 : VALUE=19'b0000000_101001101010;
      15'b010_010111000101 : VALUE=19'b0000000_101001101010;
      15'b010_010111000110 : VALUE=19'b0000000_101001101010;
      15'b010_010111000111 : VALUE=19'b0000000_101001101010;
      15'b010_010111001000 : VALUE=19'b0000000_101001101010;
      15'b010_010111001001 : VALUE=19'b0000000_101001101001;
      15'b010_010111001010 : VALUE=19'b0000000_101001101001;
      15'b010_010111001011 : VALUE=19'b0000000_101001101001;
      15'b010_010111001100 : VALUE=19'b0000000_101001101001;
      15'b010_010111001101 : VALUE=19'b0000000_101001101001;
      15'b010_010111001110 : VALUE=19'b0000000_101001101001;
      15'b010_010111001111 : VALUE=19'b0000000_101001101001;
      15'b010_010111010000 : VALUE=19'b0000000_101001101000;
      15'b010_010111010001 : VALUE=19'b0000000_101001101000;
      15'b010_010111010010 : VALUE=19'b0000000_101001101000;
      15'b010_010111010011 : VALUE=19'b0000000_101001101000;
      15'b010_010111010100 : VALUE=19'b0000000_101001101000;
      15'b010_010111010101 : VALUE=19'b0000000_101001101000;
      15'b010_010111010110 : VALUE=19'b0000000_101001101000;
      15'b010_010111010111 : VALUE=19'b0000000_101001100111;
      15'b010_010111011000 : VALUE=19'b0000000_101001100111;
      15'b010_010111011001 : VALUE=19'b0000000_101001100111;
      15'b010_010111011010 : VALUE=19'b0000000_101001100111;
      15'b010_010111011011 : VALUE=19'b0000000_101001100111;
      15'b010_010111011100 : VALUE=19'b0000000_101001100111;
      15'b010_010111011101 : VALUE=19'b0000000_101001100111;
      15'b010_010111011110 : VALUE=19'b0000000_101001100110;
      15'b010_010111011111 : VALUE=19'b0000000_101001100110;
      15'b010_010111100000 : VALUE=19'b0000000_101001100110;
      15'b010_010111100001 : VALUE=19'b0000000_101001100110;
      15'b010_010111100010 : VALUE=19'b0000000_101001100110;
      15'b010_010111100011 : VALUE=19'b0000000_101001100110;
      15'b010_010111100100 : VALUE=19'b0000000_101001100110;
      15'b010_010111100101 : VALUE=19'b0000000_101001100110;
      15'b010_010111100110 : VALUE=19'b0000000_101001100101;
      15'b010_010111100111 : VALUE=19'b0000000_101001100101;
      15'b010_010111101000 : VALUE=19'b0000000_101001100101;
      15'b010_010111101001 : VALUE=19'b0000000_101001100101;
      15'b010_010111101010 : VALUE=19'b0000000_101001100101;
      15'b010_010111101011 : VALUE=19'b0000000_101001100101;
      15'b010_010111101100 : VALUE=19'b0000000_101001100101;
      15'b010_010111101101 : VALUE=19'b0000000_101001100100;
      15'b010_010111101110 : VALUE=19'b0000000_101001100100;
      15'b010_010111101111 : VALUE=19'b0000000_101001100100;
      15'b010_010111110000 : VALUE=19'b0000000_101001100100;
      15'b010_010111110001 : VALUE=19'b0000000_101001100100;
      15'b010_010111110010 : VALUE=19'b0000000_101001100100;
      15'b010_010111110011 : VALUE=19'b0000000_101001100100;
      15'b010_010111110100 : VALUE=19'b0000000_101001100011;
      15'b010_010111110101 : VALUE=19'b0000000_101001100011;
      15'b010_010111110110 : VALUE=19'b0000000_101001100011;
      15'b010_010111110111 : VALUE=19'b0000000_101001100011;
      15'b010_010111111000 : VALUE=19'b0000000_101001100011;
      15'b010_010111111001 : VALUE=19'b0000000_101001100011;
      15'b010_010111111010 : VALUE=19'b0000000_101001100011;
      15'b010_010111111011 : VALUE=19'b0000000_101001100011;
      15'b010_010111111100 : VALUE=19'b0000000_101001100010;
      15'b010_010111111101 : VALUE=19'b0000000_101001100010;
      15'b010_010111111110 : VALUE=19'b0000000_101001100010;
      15'b010_010111111111 : VALUE=19'b0000000_101001100010;
      15'b010_011000000000 : VALUE=19'b0000000_101001100010;
      15'b010_011000000001 : VALUE=19'b0000000_101001100010;
      15'b010_011000000010 : VALUE=19'b0000000_101001100010;
      15'b010_011000000011 : VALUE=19'b0000000_101001100001;
      15'b010_011000000100 : VALUE=19'b0000000_101001100001;
      15'b010_011000000101 : VALUE=19'b0000000_101001100001;
      15'b010_011000000110 : VALUE=19'b0000000_101001100001;
      15'b010_011000000111 : VALUE=19'b0000000_101001100001;
      15'b010_011000001000 : VALUE=19'b0000000_101001100001;
      15'b010_011000001001 : VALUE=19'b0000000_101001100001;
      15'b010_011000001010 : VALUE=19'b0000000_101001100000;
      15'b010_011000001011 : VALUE=19'b0000000_101001100000;
      15'b010_011000001100 : VALUE=19'b0000000_101001100000;
      15'b010_011000001101 : VALUE=19'b0000000_101001100000;
      15'b010_011000001110 : VALUE=19'b0000000_101001100000;
      15'b010_011000001111 : VALUE=19'b0000000_101001100000;
      15'b010_011000010000 : VALUE=19'b0000000_101001100000;
      15'b010_011000010001 : VALUE=19'b0000000_101001100000;
      15'b010_011000010010 : VALUE=19'b0000000_101001011111;
      15'b010_011000010011 : VALUE=19'b0000000_101001011111;
      15'b010_011000010100 : VALUE=19'b0000000_101001011111;
      15'b010_011000010101 : VALUE=19'b0000000_101001011111;
      15'b010_011000010110 : VALUE=19'b0000000_101001011111;
      15'b010_011000010111 : VALUE=19'b0000000_101001011111;
      15'b010_011000011000 : VALUE=19'b0000000_101001011111;
      15'b010_011000011001 : VALUE=19'b0000000_101001011110;
      15'b010_011000011010 : VALUE=19'b0000000_101001011110;
      15'b010_011000011011 : VALUE=19'b0000000_101001011110;
      15'b010_011000011100 : VALUE=19'b0000000_101001011110;
      15'b010_011000011101 : VALUE=19'b0000000_101001011110;
      15'b010_011000011110 : VALUE=19'b0000000_101001011110;
      15'b010_011000011111 : VALUE=19'b0000000_101001011110;
      15'b010_011000100000 : VALUE=19'b0000000_101001011101;
      15'b010_011000100001 : VALUE=19'b0000000_101001011101;
      15'b010_011000100010 : VALUE=19'b0000000_101001011101;
      15'b010_011000100011 : VALUE=19'b0000000_101001011101;
      15'b010_011000100100 : VALUE=19'b0000000_101001011101;
      15'b010_011000100101 : VALUE=19'b0000000_101001011101;
      15'b010_011000100110 : VALUE=19'b0000000_101001011101;
      15'b010_011000100111 : VALUE=19'b0000000_101001011101;
      15'b010_011000101000 : VALUE=19'b0000000_101001011100;
      15'b010_011000101001 : VALUE=19'b0000000_101001011100;
      15'b010_011000101010 : VALUE=19'b0000000_101001011100;
      15'b010_011000101011 : VALUE=19'b0000000_101001011100;
      15'b010_011000101100 : VALUE=19'b0000000_101001011100;
      15'b010_011000101101 : VALUE=19'b0000000_101001011100;
      15'b010_011000101110 : VALUE=19'b0000000_101001011100;
      15'b010_011000101111 : VALUE=19'b0000000_101001011011;
      15'b010_011000110000 : VALUE=19'b0000000_101001011011;
      15'b010_011000110001 : VALUE=19'b0000000_101001011011;
      15'b010_011000110010 : VALUE=19'b0000000_101001011011;
      15'b010_011000110011 : VALUE=19'b0000000_101001011011;
      15'b010_011000110100 : VALUE=19'b0000000_101001011011;
      15'b010_011000110101 : VALUE=19'b0000000_101001011011;
      15'b010_011000110110 : VALUE=19'b0000000_101001011010;
      15'b010_011000110111 : VALUE=19'b0000000_101001011010;
      15'b010_011000111000 : VALUE=19'b0000000_101001011010;
      15'b010_011000111001 : VALUE=19'b0000000_101001011010;
      15'b010_011000111010 : VALUE=19'b0000000_101001011010;
      15'b010_011000111011 : VALUE=19'b0000000_101001011010;
      15'b010_011000111100 : VALUE=19'b0000000_101001011010;
      15'b010_011000111101 : VALUE=19'b0000000_101001011010;
      15'b010_011000111110 : VALUE=19'b0000000_101001011001;
      15'b010_011000111111 : VALUE=19'b0000000_101001011001;
      15'b010_011001000000 : VALUE=19'b0000000_101001011001;
      15'b010_011001000001 : VALUE=19'b0000000_101001011001;
      15'b010_011001000010 : VALUE=19'b0000000_101001011001;
      15'b010_011001000011 : VALUE=19'b0000000_101001011001;
      15'b010_011001000100 : VALUE=19'b0000000_101001011001;
      15'b010_011001000101 : VALUE=19'b0000000_101001011000;
      15'b010_011001000110 : VALUE=19'b0000000_101001011000;
      15'b010_011001000111 : VALUE=19'b0000000_101001011000;
      15'b010_011001001000 : VALUE=19'b0000000_101001011000;
      15'b010_011001001001 : VALUE=19'b0000000_101001011000;
      15'b010_011001001010 : VALUE=19'b0000000_101001011000;
      15'b010_011001001011 : VALUE=19'b0000000_101001011000;
      15'b010_011001001100 : VALUE=19'b0000000_101001011000;
      15'b010_011001001101 : VALUE=19'b0000000_101001010111;
      15'b010_011001001110 : VALUE=19'b0000000_101001010111;
      15'b010_011001001111 : VALUE=19'b0000000_101001010111;
      15'b010_011001010000 : VALUE=19'b0000000_101001010111;
      15'b010_011001010001 : VALUE=19'b0000000_101001010111;
      15'b010_011001010010 : VALUE=19'b0000000_101001010111;
      15'b010_011001010011 : VALUE=19'b0000000_101001010111;
      15'b010_011001010100 : VALUE=19'b0000000_101001010110;
      15'b010_011001010101 : VALUE=19'b0000000_101001010110;
      15'b010_011001010110 : VALUE=19'b0000000_101001010110;
      15'b010_011001010111 : VALUE=19'b0000000_101001010110;
      15'b010_011001011000 : VALUE=19'b0000000_101001010110;
      15'b010_011001011001 : VALUE=19'b0000000_101001010110;
      15'b010_011001011010 : VALUE=19'b0000000_101001010110;
      15'b010_011001011011 : VALUE=19'b0000000_101001010101;
      15'b010_011001011100 : VALUE=19'b0000000_101001010101;
      15'b010_011001011101 : VALUE=19'b0000000_101001010101;
      15'b010_011001011110 : VALUE=19'b0000000_101001010101;
      15'b010_011001011111 : VALUE=19'b0000000_101001010101;
      15'b010_011001100000 : VALUE=19'b0000000_101001010101;
      15'b010_011001100001 : VALUE=19'b0000000_101001010101;
      15'b010_011001100010 : VALUE=19'b0000000_101001010101;
      15'b010_011001100011 : VALUE=19'b0000000_101001010100;
      15'b010_011001100100 : VALUE=19'b0000000_101001010100;
      15'b010_011001100101 : VALUE=19'b0000000_101001010100;
      15'b010_011001100110 : VALUE=19'b0000000_101001010100;
      15'b010_011001100111 : VALUE=19'b0000000_101001010100;
      15'b010_011001101000 : VALUE=19'b0000000_101001010100;
      15'b010_011001101001 : VALUE=19'b0000000_101001010100;
      15'b010_011001101010 : VALUE=19'b0000000_101001010011;
      15'b010_011001101011 : VALUE=19'b0000000_101001010011;
      15'b010_011001101100 : VALUE=19'b0000000_101001010011;
      15'b010_011001101101 : VALUE=19'b0000000_101001010011;
      15'b010_011001101110 : VALUE=19'b0000000_101001010011;
      15'b010_011001101111 : VALUE=19'b0000000_101001010011;
      15'b010_011001110000 : VALUE=19'b0000000_101001010011;
      15'b010_011001110001 : VALUE=19'b0000000_101001010011;
      15'b010_011001110010 : VALUE=19'b0000000_101001010010;
      15'b010_011001110011 : VALUE=19'b0000000_101001010010;
      15'b010_011001110100 : VALUE=19'b0000000_101001010010;
      15'b010_011001110101 : VALUE=19'b0000000_101001010010;
      15'b010_011001110110 : VALUE=19'b0000000_101001010010;
      15'b010_011001110111 : VALUE=19'b0000000_101001010010;
      15'b010_011001111000 : VALUE=19'b0000000_101001010010;
      15'b010_011001111001 : VALUE=19'b0000000_101001010001;
      15'b010_011001111010 : VALUE=19'b0000000_101001010001;
      15'b010_011001111011 : VALUE=19'b0000000_101001010001;
      15'b010_011001111100 : VALUE=19'b0000000_101001010001;
      15'b010_011001111101 : VALUE=19'b0000000_101001010001;
      15'b010_011001111110 : VALUE=19'b0000000_101001010001;
      15'b010_011001111111 : VALUE=19'b0000000_101001010001;
      15'b010_011010000000 : VALUE=19'b0000000_101001010001;
      15'b010_011010000001 : VALUE=19'b0000000_101001010000;
      15'b010_011010000010 : VALUE=19'b0000000_101001010000;
      15'b010_011010000011 : VALUE=19'b0000000_101001010000;
      15'b010_011010000100 : VALUE=19'b0000000_101001010000;
      15'b010_011010000101 : VALUE=19'b0000000_101001010000;
      15'b010_011010000110 : VALUE=19'b0000000_101001010000;
      15'b010_011010000111 : VALUE=19'b0000000_101001010000;
      15'b010_011010001000 : VALUE=19'b0000000_101001001111;
      15'b010_011010001001 : VALUE=19'b0000000_101001001111;
      15'b010_011010001010 : VALUE=19'b0000000_101001001111;
      15'b010_011010001011 : VALUE=19'b0000000_101001001111;
      15'b010_011010001100 : VALUE=19'b0000000_101001001111;
      15'b010_011010001101 : VALUE=19'b0000000_101001001111;
      15'b010_011010001110 : VALUE=19'b0000000_101001001111;
      15'b010_011010001111 : VALUE=19'b0000000_101001001111;
      15'b010_011010010000 : VALUE=19'b0000000_101001001110;
      15'b010_011010010001 : VALUE=19'b0000000_101001001110;
      15'b010_011010010010 : VALUE=19'b0000000_101001001110;
      15'b010_011010010011 : VALUE=19'b0000000_101001001110;
      15'b010_011010010100 : VALUE=19'b0000000_101001001110;
      15'b010_011010010101 : VALUE=19'b0000000_101001001110;
      15'b010_011010010110 : VALUE=19'b0000000_101001001110;
      15'b010_011010010111 : VALUE=19'b0000000_101001001101;
      15'b010_011010011000 : VALUE=19'b0000000_101001001101;
      15'b010_011010011001 : VALUE=19'b0000000_101001001101;
      15'b010_011010011010 : VALUE=19'b0000000_101001001101;
      15'b010_011010011011 : VALUE=19'b0000000_101001001101;
      15'b010_011010011100 : VALUE=19'b0000000_101001001101;
      15'b010_011010011101 : VALUE=19'b0000000_101001001101;
      15'b010_011010011110 : VALUE=19'b0000000_101001001101;
      15'b010_011010011111 : VALUE=19'b0000000_101001001100;
      15'b010_011010100000 : VALUE=19'b0000000_101001001100;
      15'b010_011010100001 : VALUE=19'b0000000_101001001100;
      15'b010_011010100010 : VALUE=19'b0000000_101001001100;
      15'b010_011010100011 : VALUE=19'b0000000_101001001100;
      15'b010_011010100100 : VALUE=19'b0000000_101001001100;
      15'b010_011010100101 : VALUE=19'b0000000_101001001100;
      15'b010_011010100110 : VALUE=19'b0000000_101001001011;
      15'b010_011010100111 : VALUE=19'b0000000_101001001011;
      15'b010_011010101000 : VALUE=19'b0000000_101001001011;
      15'b010_011010101001 : VALUE=19'b0000000_101001001011;
      15'b010_011010101010 : VALUE=19'b0000000_101001001011;
      15'b010_011010101011 : VALUE=19'b0000000_101001001011;
      15'b010_011010101100 : VALUE=19'b0000000_101001001011;
      15'b010_011010101101 : VALUE=19'b0000000_101001001011;
      15'b010_011010101110 : VALUE=19'b0000000_101001001010;
      15'b010_011010101111 : VALUE=19'b0000000_101001001010;
      15'b010_011010110000 : VALUE=19'b0000000_101001001010;
      15'b010_011010110001 : VALUE=19'b0000000_101001001010;
      15'b010_011010110010 : VALUE=19'b0000000_101001001010;
      15'b010_011010110011 : VALUE=19'b0000000_101001001010;
      15'b010_011010110100 : VALUE=19'b0000000_101001001010;
      15'b010_011010110101 : VALUE=19'b0000000_101001001001;
      15'b010_011010110110 : VALUE=19'b0000000_101001001001;
      15'b010_011010110111 : VALUE=19'b0000000_101001001001;
      15'b010_011010111000 : VALUE=19'b0000000_101001001001;
      15'b010_011010111001 : VALUE=19'b0000000_101001001001;
      15'b010_011010111010 : VALUE=19'b0000000_101001001001;
      15'b010_011010111011 : VALUE=19'b0000000_101001001001;
      15'b010_011010111100 : VALUE=19'b0000000_101001001001;
      15'b010_011010111101 : VALUE=19'b0000000_101001001000;
      15'b010_011010111110 : VALUE=19'b0000000_101001001000;
      15'b010_011010111111 : VALUE=19'b0000000_101001001000;
      15'b010_011011000000 : VALUE=19'b0000000_101001001000;
      15'b010_011011000001 : VALUE=19'b0000000_101001001000;
      15'b010_011011000010 : VALUE=19'b0000000_101001001000;
      15'b010_011011000011 : VALUE=19'b0000000_101001001000;
      15'b010_011011000100 : VALUE=19'b0000000_101001000111;
      15'b010_011011000101 : VALUE=19'b0000000_101001000111;
      15'b010_011011000110 : VALUE=19'b0000000_101001000111;
      15'b010_011011000111 : VALUE=19'b0000000_101001000111;
      15'b010_011011001000 : VALUE=19'b0000000_101001000111;
      15'b010_011011001001 : VALUE=19'b0000000_101001000111;
      15'b010_011011001010 : VALUE=19'b0000000_101001000111;
      15'b010_011011001011 : VALUE=19'b0000000_101001000111;
      15'b010_011011001100 : VALUE=19'b0000000_101001000110;
      15'b010_011011001101 : VALUE=19'b0000000_101001000110;
      15'b010_011011001110 : VALUE=19'b0000000_101001000110;
      15'b010_011011001111 : VALUE=19'b0000000_101001000110;
      15'b010_011011010000 : VALUE=19'b0000000_101001000110;
      15'b010_011011010001 : VALUE=19'b0000000_101001000110;
      15'b010_011011010010 : VALUE=19'b0000000_101001000110;
      15'b010_011011010011 : VALUE=19'b0000000_101001000101;
      15'b010_011011010100 : VALUE=19'b0000000_101001000101;
      15'b010_011011010101 : VALUE=19'b0000000_101001000101;
      15'b010_011011010110 : VALUE=19'b0000000_101001000101;
      15'b010_011011010111 : VALUE=19'b0000000_101001000101;
      15'b010_011011011000 : VALUE=19'b0000000_101001000101;
      15'b010_011011011001 : VALUE=19'b0000000_101001000101;
      15'b010_011011011010 : VALUE=19'b0000000_101001000101;
      15'b010_011011011011 : VALUE=19'b0000000_101001000100;
      15'b010_011011011100 : VALUE=19'b0000000_101001000100;
      15'b010_011011011101 : VALUE=19'b0000000_101001000100;
      15'b010_011011011110 : VALUE=19'b0000000_101001000100;
      15'b010_011011011111 : VALUE=19'b0000000_101001000100;
      15'b010_011011100000 : VALUE=19'b0000000_101001000100;
      15'b010_011011100001 : VALUE=19'b0000000_101001000100;
      15'b010_011011100010 : VALUE=19'b0000000_101001000011;
      15'b010_011011100011 : VALUE=19'b0000000_101001000011;
      15'b010_011011100100 : VALUE=19'b0000000_101001000011;
      15'b010_011011100101 : VALUE=19'b0000000_101001000011;
      15'b010_011011100110 : VALUE=19'b0000000_101001000011;
      15'b010_011011100111 : VALUE=19'b0000000_101001000011;
      15'b010_011011101000 : VALUE=19'b0000000_101001000011;
      15'b010_011011101001 : VALUE=19'b0000000_101001000011;
      15'b010_011011101010 : VALUE=19'b0000000_101001000010;
      15'b010_011011101011 : VALUE=19'b0000000_101001000010;
      15'b010_011011101100 : VALUE=19'b0000000_101001000010;
      15'b010_011011101101 : VALUE=19'b0000000_101001000010;
      15'b010_011011101110 : VALUE=19'b0000000_101001000010;
      15'b010_011011101111 : VALUE=19'b0000000_101001000010;
      15'b010_011011110000 : VALUE=19'b0000000_101001000010;
      15'b010_011011110001 : VALUE=19'b0000000_101001000010;
      15'b010_011011110010 : VALUE=19'b0000000_101001000001;
      15'b010_011011110011 : VALUE=19'b0000000_101001000001;
      15'b010_011011110100 : VALUE=19'b0000000_101001000001;
      15'b010_011011110101 : VALUE=19'b0000000_101001000001;
      15'b010_011011110110 : VALUE=19'b0000000_101001000001;
      15'b010_011011110111 : VALUE=19'b0000000_101001000001;
      15'b010_011011111000 : VALUE=19'b0000000_101001000001;
      15'b010_011011111001 : VALUE=19'b0000000_101001000000;
      15'b010_011011111010 : VALUE=19'b0000000_101001000000;
      15'b010_011011111011 : VALUE=19'b0000000_101001000000;
      15'b010_011011111100 : VALUE=19'b0000000_101001000000;
      15'b010_011011111101 : VALUE=19'b0000000_101001000000;
      15'b010_011011111110 : VALUE=19'b0000000_101001000000;
      15'b010_011011111111 : VALUE=19'b0000000_101001000000;
      15'b010_011100000000 : VALUE=19'b0000000_101001000000;
      15'b010_011100000001 : VALUE=19'b0000000_101000111111;
      15'b010_011100000010 : VALUE=19'b0000000_101000111111;
      15'b010_011100000011 : VALUE=19'b0000000_101000111111;
      15'b010_011100000100 : VALUE=19'b0000000_101000111111;
      15'b010_011100000101 : VALUE=19'b0000000_101000111111;
      15'b010_011100000110 : VALUE=19'b0000000_101000111111;
      15'b010_011100000111 : VALUE=19'b0000000_101000111111;
      15'b010_011100001000 : VALUE=19'b0000000_101000111110;
      15'b010_011100001001 : VALUE=19'b0000000_101000111110;
      15'b010_011100001010 : VALUE=19'b0000000_101000111110;
      15'b010_011100001011 : VALUE=19'b0000000_101000111110;
      15'b010_011100001100 : VALUE=19'b0000000_101000111110;
      15'b010_011100001101 : VALUE=19'b0000000_101000111110;
      15'b010_011100001110 : VALUE=19'b0000000_101000111110;
      15'b010_011100001111 : VALUE=19'b0000000_101000111110;
      15'b010_011100010000 : VALUE=19'b0000000_101000111101;
      15'b010_011100010001 : VALUE=19'b0000000_101000111101;
      15'b010_011100010010 : VALUE=19'b0000000_101000111101;
      15'b010_011100010011 : VALUE=19'b0000000_101000111101;
      15'b010_011100010100 : VALUE=19'b0000000_101000111101;
      15'b010_011100010101 : VALUE=19'b0000000_101000111101;
      15'b010_011100010110 : VALUE=19'b0000000_101000111101;
      15'b010_011100010111 : VALUE=19'b0000000_101000111101;
      15'b010_011100011000 : VALUE=19'b0000000_101000111100;
      15'b010_011100011001 : VALUE=19'b0000000_101000111100;
      15'b010_011100011010 : VALUE=19'b0000000_101000111100;
      15'b010_011100011011 : VALUE=19'b0000000_101000111100;
      15'b010_011100011100 : VALUE=19'b0000000_101000111100;
      15'b010_011100011101 : VALUE=19'b0000000_101000111100;
      15'b010_011100011110 : VALUE=19'b0000000_101000111100;
      15'b010_011100011111 : VALUE=19'b0000000_101000111011;
      15'b010_011100100000 : VALUE=19'b0000000_101000111011;
      15'b010_011100100001 : VALUE=19'b0000000_101000111011;
      15'b010_011100100010 : VALUE=19'b0000000_101000111011;
      15'b010_011100100011 : VALUE=19'b0000000_101000111011;
      15'b010_011100100100 : VALUE=19'b0000000_101000111011;
      15'b010_011100100101 : VALUE=19'b0000000_101000111011;
      15'b010_011100100110 : VALUE=19'b0000000_101000111011;
      15'b010_011100100111 : VALUE=19'b0000000_101000111010;
      15'b010_011100101000 : VALUE=19'b0000000_101000111010;
      15'b010_011100101001 : VALUE=19'b0000000_101000111010;
      15'b010_011100101010 : VALUE=19'b0000000_101000111010;
      15'b010_011100101011 : VALUE=19'b0000000_101000111010;
      15'b010_011100101100 : VALUE=19'b0000000_101000111010;
      15'b010_011100101101 : VALUE=19'b0000000_101000111010;
      15'b010_011100101110 : VALUE=19'b0000000_101000111010;
      15'b010_011100101111 : VALUE=19'b0000000_101000111001;
      15'b010_011100110000 : VALUE=19'b0000000_101000111001;
      15'b010_011100110001 : VALUE=19'b0000000_101000111001;
      15'b010_011100110010 : VALUE=19'b0000000_101000111001;
      15'b010_011100110011 : VALUE=19'b0000000_101000111001;
      15'b010_011100110100 : VALUE=19'b0000000_101000111001;
      15'b010_011100110101 : VALUE=19'b0000000_101000111001;
      15'b010_011100110110 : VALUE=19'b0000000_101000111000;
      15'b010_011100110111 : VALUE=19'b0000000_101000111000;
      15'b010_011100111000 : VALUE=19'b0000000_101000111000;
      15'b010_011100111001 : VALUE=19'b0000000_101000111000;
      15'b010_011100111010 : VALUE=19'b0000000_101000111000;
      15'b010_011100111011 : VALUE=19'b0000000_101000111000;
      15'b010_011100111100 : VALUE=19'b0000000_101000111000;
      15'b010_011100111101 : VALUE=19'b0000000_101000111000;
      15'b010_011100111110 : VALUE=19'b0000000_101000110111;
      15'b010_011100111111 : VALUE=19'b0000000_101000110111;
      15'b010_011101000000 : VALUE=19'b0000000_101000110111;
      15'b010_011101000001 : VALUE=19'b0000000_101000110111;
      15'b010_011101000010 : VALUE=19'b0000000_101000110111;
      15'b010_011101000011 : VALUE=19'b0000000_101000110111;
      15'b010_011101000100 : VALUE=19'b0000000_101000110111;
      15'b010_011101000101 : VALUE=19'b0000000_101000110111;
      15'b010_011101000110 : VALUE=19'b0000000_101000110110;
      15'b010_011101000111 : VALUE=19'b0000000_101000110110;
      15'b010_011101001000 : VALUE=19'b0000000_101000110110;
      15'b010_011101001001 : VALUE=19'b0000000_101000110110;
      15'b010_011101001010 : VALUE=19'b0000000_101000110110;
      15'b010_011101001011 : VALUE=19'b0000000_101000110110;
      15'b010_011101001100 : VALUE=19'b0000000_101000110110;
      15'b010_011101001101 : VALUE=19'b0000000_101000110101;
      15'b010_011101001110 : VALUE=19'b0000000_101000110101;
      15'b010_011101001111 : VALUE=19'b0000000_101000110101;
      15'b010_011101010000 : VALUE=19'b0000000_101000110101;
      15'b010_011101010001 : VALUE=19'b0000000_101000110101;
      15'b010_011101010010 : VALUE=19'b0000000_101000110101;
      15'b010_011101010011 : VALUE=19'b0000000_101000110101;
      15'b010_011101010100 : VALUE=19'b0000000_101000110101;
      15'b010_011101010101 : VALUE=19'b0000000_101000110100;
      15'b010_011101010110 : VALUE=19'b0000000_101000110100;
      15'b010_011101010111 : VALUE=19'b0000000_101000110100;
      15'b010_011101011000 : VALUE=19'b0000000_101000110100;
      15'b010_011101011001 : VALUE=19'b0000000_101000110100;
      15'b010_011101011010 : VALUE=19'b0000000_101000110100;
      15'b010_011101011011 : VALUE=19'b0000000_101000110100;
      15'b010_011101011100 : VALUE=19'b0000000_101000110100;
      15'b010_011101011101 : VALUE=19'b0000000_101000110011;
      15'b010_011101011110 : VALUE=19'b0000000_101000110011;
      15'b010_011101011111 : VALUE=19'b0000000_101000110011;
      15'b010_011101100000 : VALUE=19'b0000000_101000110011;
      15'b010_011101100001 : VALUE=19'b0000000_101000110011;
      15'b010_011101100010 : VALUE=19'b0000000_101000110011;
      15'b010_011101100011 : VALUE=19'b0000000_101000110011;
      15'b010_011101100100 : VALUE=19'b0000000_101000110010;
      15'b010_011101100101 : VALUE=19'b0000000_101000110010;
      15'b010_011101100110 : VALUE=19'b0000000_101000110010;
      15'b010_011101100111 : VALUE=19'b0000000_101000110010;
      15'b010_011101101000 : VALUE=19'b0000000_101000110010;
      15'b010_011101101001 : VALUE=19'b0000000_101000110010;
      15'b010_011101101010 : VALUE=19'b0000000_101000110010;
      15'b010_011101101011 : VALUE=19'b0000000_101000110010;
      15'b010_011101101100 : VALUE=19'b0000000_101000110001;
      15'b010_011101101101 : VALUE=19'b0000000_101000110001;
      15'b010_011101101110 : VALUE=19'b0000000_101000110001;
      15'b010_011101101111 : VALUE=19'b0000000_101000110001;
      15'b010_011101110000 : VALUE=19'b0000000_101000110001;
      15'b010_011101110001 : VALUE=19'b0000000_101000110001;
      15'b010_011101110010 : VALUE=19'b0000000_101000110001;
      15'b010_011101110011 : VALUE=19'b0000000_101000110001;
      15'b010_011101110100 : VALUE=19'b0000000_101000110000;
      15'b010_011101110101 : VALUE=19'b0000000_101000110000;
      15'b010_011101110110 : VALUE=19'b0000000_101000110000;
      15'b010_011101110111 : VALUE=19'b0000000_101000110000;
      15'b010_011101111000 : VALUE=19'b0000000_101000110000;
      15'b010_011101111001 : VALUE=19'b0000000_101000110000;
      15'b010_011101111010 : VALUE=19'b0000000_101000110000;
      15'b010_011101111011 : VALUE=19'b0000000_101000110000;
      15'b010_011101111100 : VALUE=19'b0000000_101000101111;
      15'b010_011101111101 : VALUE=19'b0000000_101000101111;
      15'b010_011101111110 : VALUE=19'b0000000_101000101111;
      15'b010_011101111111 : VALUE=19'b0000000_101000101111;
      15'b010_011110000000 : VALUE=19'b0000000_101000101111;
      15'b010_011110000001 : VALUE=19'b0000000_101000101111;
      15'b010_011110000010 : VALUE=19'b0000000_101000101111;
      15'b010_011110000011 : VALUE=19'b0000000_101000101110;
      15'b010_011110000100 : VALUE=19'b0000000_101000101110;
      15'b010_011110000101 : VALUE=19'b0000000_101000101110;
      15'b010_011110000110 : VALUE=19'b0000000_101000101110;
      15'b010_011110000111 : VALUE=19'b0000000_101000101110;
      15'b010_011110001000 : VALUE=19'b0000000_101000101110;
      15'b010_011110001001 : VALUE=19'b0000000_101000101110;
      15'b010_011110001010 : VALUE=19'b0000000_101000101110;
      15'b010_011110001011 : VALUE=19'b0000000_101000101101;
      15'b010_011110001100 : VALUE=19'b0000000_101000101101;
      15'b010_011110001101 : VALUE=19'b0000000_101000101101;
      15'b010_011110001110 : VALUE=19'b0000000_101000101101;
      15'b010_011110001111 : VALUE=19'b0000000_101000101101;
      15'b010_011110010000 : VALUE=19'b0000000_101000101101;
      15'b010_011110010001 : VALUE=19'b0000000_101000101101;
      15'b010_011110010010 : VALUE=19'b0000000_101000101101;
      15'b010_011110010011 : VALUE=19'b0000000_101000101100;
      15'b010_011110010100 : VALUE=19'b0000000_101000101100;
      15'b010_011110010101 : VALUE=19'b0000000_101000101100;
      15'b010_011110010110 : VALUE=19'b0000000_101000101100;
      15'b010_011110010111 : VALUE=19'b0000000_101000101100;
      15'b010_011110011000 : VALUE=19'b0000000_101000101100;
      15'b010_011110011001 : VALUE=19'b0000000_101000101100;
      15'b010_011110011010 : VALUE=19'b0000000_101000101100;
      15'b010_011110011011 : VALUE=19'b0000000_101000101011;
      15'b010_011110011100 : VALUE=19'b0000000_101000101011;
      15'b010_011110011101 : VALUE=19'b0000000_101000101011;
      15'b010_011110011110 : VALUE=19'b0000000_101000101011;
      15'b010_011110011111 : VALUE=19'b0000000_101000101011;
      15'b010_011110100000 : VALUE=19'b0000000_101000101011;
      15'b010_011110100001 : VALUE=19'b0000000_101000101011;
      15'b010_011110100010 : VALUE=19'b0000000_101000101011;
      15'b010_011110100011 : VALUE=19'b0000000_101000101010;
      15'b010_011110100100 : VALUE=19'b0000000_101000101010;
      15'b010_011110100101 : VALUE=19'b0000000_101000101010;
      15'b010_011110100110 : VALUE=19'b0000000_101000101010;
      15'b010_011110100111 : VALUE=19'b0000000_101000101010;
      15'b010_011110101000 : VALUE=19'b0000000_101000101010;
      15'b010_011110101001 : VALUE=19'b0000000_101000101010;
      15'b010_011110101010 : VALUE=19'b0000000_101000101001;
      15'b010_011110101011 : VALUE=19'b0000000_101000101001;
      15'b010_011110101100 : VALUE=19'b0000000_101000101001;
      15'b010_011110101101 : VALUE=19'b0000000_101000101001;
      15'b010_011110101110 : VALUE=19'b0000000_101000101001;
      15'b010_011110101111 : VALUE=19'b0000000_101000101001;
      15'b010_011110110000 : VALUE=19'b0000000_101000101001;
      15'b010_011110110001 : VALUE=19'b0000000_101000101001;
      15'b010_011110110010 : VALUE=19'b0000000_101000101000;
      15'b010_011110110011 : VALUE=19'b0000000_101000101000;
      15'b010_011110110100 : VALUE=19'b0000000_101000101000;
      15'b010_011110110101 : VALUE=19'b0000000_101000101000;
      15'b010_011110110110 : VALUE=19'b0000000_101000101000;
      15'b010_011110110111 : VALUE=19'b0000000_101000101000;
      15'b010_011110111000 : VALUE=19'b0000000_101000101000;
      15'b010_011110111001 : VALUE=19'b0000000_101000101000;
      15'b010_011110111010 : VALUE=19'b0000000_101000100111;
      15'b010_011110111011 : VALUE=19'b0000000_101000100111;
      15'b010_011110111100 : VALUE=19'b0000000_101000100111;
      15'b010_011110111101 : VALUE=19'b0000000_101000100111;
      15'b010_011110111110 : VALUE=19'b0000000_101000100111;
      15'b010_011110111111 : VALUE=19'b0000000_101000100111;
      15'b010_011111000000 : VALUE=19'b0000000_101000100111;
      15'b010_011111000001 : VALUE=19'b0000000_101000100111;
      15'b010_011111000010 : VALUE=19'b0000000_101000100110;
      15'b010_011111000011 : VALUE=19'b0000000_101000100110;
      15'b010_011111000100 : VALUE=19'b0000000_101000100110;
      15'b010_011111000101 : VALUE=19'b0000000_101000100110;
      15'b010_011111000110 : VALUE=19'b0000000_101000100110;
      15'b010_011111000111 : VALUE=19'b0000000_101000100110;
      15'b010_011111001000 : VALUE=19'b0000000_101000100110;
      15'b010_011111001001 : VALUE=19'b0000000_101000100110;
      15'b010_011111001010 : VALUE=19'b0000000_101000100101;
      15'b010_011111001011 : VALUE=19'b0000000_101000100101;
      15'b010_011111001100 : VALUE=19'b0000000_101000100101;
      15'b010_011111001101 : VALUE=19'b0000000_101000100101;
      15'b010_011111001110 : VALUE=19'b0000000_101000100101;
      15'b010_011111001111 : VALUE=19'b0000000_101000100101;
      15'b010_011111010000 : VALUE=19'b0000000_101000100101;
      15'b010_011111010001 : VALUE=19'b0000000_101000100101;
      15'b010_011111010010 : VALUE=19'b0000000_101000100100;
      15'b010_011111010011 : VALUE=19'b0000000_101000100100;
      15'b010_011111010100 : VALUE=19'b0000000_101000100100;
      15'b010_011111010101 : VALUE=19'b0000000_101000100100;
      15'b010_011111010110 : VALUE=19'b0000000_101000100100;
      15'b010_011111010111 : VALUE=19'b0000000_101000100100;
      15'b010_011111011000 : VALUE=19'b0000000_101000100100;
      15'b010_011111011001 : VALUE=19'b0000000_101000100011;
      15'b010_011111011010 : VALUE=19'b0000000_101000100011;
      15'b010_011111011011 : VALUE=19'b0000000_101000100011;
      15'b010_011111011100 : VALUE=19'b0000000_101000100011;
      15'b010_011111011101 : VALUE=19'b0000000_101000100011;
      15'b010_011111011110 : VALUE=19'b0000000_101000100011;
      15'b010_011111011111 : VALUE=19'b0000000_101000100011;
      15'b010_011111100000 : VALUE=19'b0000000_101000100011;
      15'b010_011111100001 : VALUE=19'b0000000_101000100010;
      15'b010_011111100010 : VALUE=19'b0000000_101000100010;
      15'b010_011111100011 : VALUE=19'b0000000_101000100010;
      15'b010_011111100100 : VALUE=19'b0000000_101000100010;
      15'b010_011111100101 : VALUE=19'b0000000_101000100010;
      15'b010_011111100110 : VALUE=19'b0000000_101000100010;
      15'b010_011111100111 : VALUE=19'b0000000_101000100010;
      15'b010_011111101000 : VALUE=19'b0000000_101000100010;
      15'b010_011111101001 : VALUE=19'b0000000_101000100001;
      15'b010_011111101010 : VALUE=19'b0000000_101000100001;
      15'b010_011111101011 : VALUE=19'b0000000_101000100001;
      15'b010_011111101100 : VALUE=19'b0000000_101000100001;
      15'b010_011111101101 : VALUE=19'b0000000_101000100001;
      15'b010_011111101110 : VALUE=19'b0000000_101000100001;
      15'b010_011111101111 : VALUE=19'b0000000_101000100001;
      15'b010_011111110000 : VALUE=19'b0000000_101000100001;
      15'b010_011111110001 : VALUE=19'b0000000_101000100000;
      15'b010_011111110010 : VALUE=19'b0000000_101000100000;
      15'b010_011111110011 : VALUE=19'b0000000_101000100000;
      15'b010_011111110100 : VALUE=19'b0000000_101000100000;
      15'b010_011111110101 : VALUE=19'b0000000_101000100000;
      15'b010_011111110110 : VALUE=19'b0000000_101000100000;
      15'b010_011111110111 : VALUE=19'b0000000_101000100000;
      15'b010_011111111000 : VALUE=19'b0000000_101000100000;
      15'b010_011111111001 : VALUE=19'b0000000_101000011111;
      15'b010_011111111010 : VALUE=19'b0000000_101000011111;
      15'b010_011111111011 : VALUE=19'b0000000_101000011111;
      15'b010_011111111100 : VALUE=19'b0000000_101000011111;
      15'b010_011111111101 : VALUE=19'b0000000_101000011111;
      15'b010_011111111110 : VALUE=19'b0000000_101000011111;
      15'b010_011111111111 : VALUE=19'b0000000_101000011111;
      15'b010_100000000000 : VALUE=19'b0000000_101000011111;
      15'b010_100000000001 : VALUE=19'b0000000_101000011110;
      15'b010_100000000010 : VALUE=19'b0000000_101000011110;
      15'b010_100000000011 : VALUE=19'b0000000_101000011110;
      15'b010_100000000100 : VALUE=19'b0000000_101000011110;
      15'b010_100000000101 : VALUE=19'b0000000_101000011110;
      15'b010_100000000110 : VALUE=19'b0000000_101000011110;
      15'b010_100000000111 : VALUE=19'b0000000_101000011110;
      15'b010_100000001000 : VALUE=19'b0000000_101000011110;
      15'b010_100000001001 : VALUE=19'b0000000_101000011101;
      15'b010_100000001010 : VALUE=19'b0000000_101000011101;
      15'b010_100000001011 : VALUE=19'b0000000_101000011101;
      15'b010_100000001100 : VALUE=19'b0000000_101000011101;
      15'b010_100000001101 : VALUE=19'b0000000_101000011101;
      15'b010_100000001110 : VALUE=19'b0000000_101000011101;
      15'b010_100000001111 : VALUE=19'b0000000_101000011101;
      15'b010_100000010000 : VALUE=19'b0000000_101000011101;
      15'b010_100000010001 : VALUE=19'b0000000_101000011100;
      15'b010_100000010010 : VALUE=19'b0000000_101000011100;
      15'b010_100000010011 : VALUE=19'b0000000_101000011100;
      15'b010_100000010100 : VALUE=19'b0000000_101000011100;
      15'b010_100000010101 : VALUE=19'b0000000_101000011100;
      15'b010_100000010110 : VALUE=19'b0000000_101000011100;
      15'b010_100000010111 : VALUE=19'b0000000_101000011100;
      15'b010_100000011000 : VALUE=19'b0000000_101000011100;
      15'b010_100000011001 : VALUE=19'b0000000_101000011011;
      15'b010_100000011010 : VALUE=19'b0000000_101000011011;
      15'b010_100000011011 : VALUE=19'b0000000_101000011011;
      15'b010_100000011100 : VALUE=19'b0000000_101000011011;
      15'b010_100000011101 : VALUE=19'b0000000_101000011011;
      15'b010_100000011110 : VALUE=19'b0000000_101000011011;
      15'b010_100000011111 : VALUE=19'b0000000_101000011011;
      15'b010_100000100000 : VALUE=19'b0000000_101000011010;
      15'b010_100000100001 : VALUE=19'b0000000_101000011010;
      15'b010_100000100010 : VALUE=19'b0000000_101000011010;
      15'b010_100000100011 : VALUE=19'b0000000_101000011010;
      15'b010_100000100100 : VALUE=19'b0000000_101000011010;
      15'b010_100000100101 : VALUE=19'b0000000_101000011010;
      15'b010_100000100110 : VALUE=19'b0000000_101000011010;
      15'b010_100000100111 : VALUE=19'b0000000_101000011010;
      15'b010_100000101000 : VALUE=19'b0000000_101000011001;
      15'b010_100000101001 : VALUE=19'b0000000_101000011001;
      15'b010_100000101010 : VALUE=19'b0000000_101000011001;
      15'b010_100000101011 : VALUE=19'b0000000_101000011001;
      15'b010_100000101100 : VALUE=19'b0000000_101000011001;
      15'b010_100000101101 : VALUE=19'b0000000_101000011001;
      15'b010_100000101110 : VALUE=19'b0000000_101000011001;
      15'b010_100000101111 : VALUE=19'b0000000_101000011001;
      15'b010_100000110000 : VALUE=19'b0000000_101000011000;
      15'b010_100000110001 : VALUE=19'b0000000_101000011000;
      15'b010_100000110010 : VALUE=19'b0000000_101000011000;
      15'b010_100000110011 : VALUE=19'b0000000_101000011000;
      15'b010_100000110100 : VALUE=19'b0000000_101000011000;
      15'b010_100000110101 : VALUE=19'b0000000_101000011000;
      15'b010_100000110110 : VALUE=19'b0000000_101000011000;
      15'b010_100000110111 : VALUE=19'b0000000_101000011000;
      15'b010_100000111000 : VALUE=19'b0000000_101000010111;
      15'b010_100000111001 : VALUE=19'b0000000_101000010111;
      15'b010_100000111010 : VALUE=19'b0000000_101000010111;
      15'b010_100000111011 : VALUE=19'b0000000_101000010111;
      15'b010_100000111100 : VALUE=19'b0000000_101000010111;
      15'b010_100000111101 : VALUE=19'b0000000_101000010111;
      15'b010_100000111110 : VALUE=19'b0000000_101000010111;
      15'b010_100000111111 : VALUE=19'b0000000_101000010111;
      15'b010_100001000000 : VALUE=19'b0000000_101000010110;
      15'b010_100001000001 : VALUE=19'b0000000_101000010110;
      15'b010_100001000010 : VALUE=19'b0000000_101000010110;
      15'b010_100001000011 : VALUE=19'b0000000_101000010110;
      15'b010_100001000100 : VALUE=19'b0000000_101000010110;
      15'b010_100001000101 : VALUE=19'b0000000_101000010110;
      15'b010_100001000110 : VALUE=19'b0000000_101000010110;
      15'b010_100001000111 : VALUE=19'b0000000_101000010110;
      15'b010_100001001000 : VALUE=19'b0000000_101000010101;
      15'b010_100001001001 : VALUE=19'b0000000_101000010101;
      15'b010_100001001010 : VALUE=19'b0000000_101000010101;
      15'b010_100001001011 : VALUE=19'b0000000_101000010101;
      15'b010_100001001100 : VALUE=19'b0000000_101000010101;
      15'b010_100001001101 : VALUE=19'b0000000_101000010101;
      15'b010_100001001110 : VALUE=19'b0000000_101000010101;
      15'b010_100001001111 : VALUE=19'b0000000_101000010101;
      15'b010_100001010000 : VALUE=19'b0000000_101000010100;
      15'b010_100001010001 : VALUE=19'b0000000_101000010100;
      15'b010_100001010010 : VALUE=19'b0000000_101000010100;
      15'b010_100001010011 : VALUE=19'b0000000_101000010100;
      15'b010_100001010100 : VALUE=19'b0000000_101000010100;
      15'b010_100001010101 : VALUE=19'b0000000_101000010100;
      15'b010_100001010110 : VALUE=19'b0000000_101000010100;
      15'b010_100001010111 : VALUE=19'b0000000_101000010100;
      15'b010_100001011000 : VALUE=19'b0000000_101000010011;
      15'b010_100001011001 : VALUE=19'b0000000_101000010011;
      15'b010_100001011010 : VALUE=19'b0000000_101000010011;
      15'b010_100001011011 : VALUE=19'b0000000_101000010011;
      15'b010_100001011100 : VALUE=19'b0000000_101000010011;
      15'b010_100001011101 : VALUE=19'b0000000_101000010011;
      15'b010_100001011110 : VALUE=19'b0000000_101000010011;
      15'b010_100001011111 : VALUE=19'b0000000_101000010011;
      15'b010_100001100000 : VALUE=19'b0000000_101000010010;
      15'b010_100001100001 : VALUE=19'b0000000_101000010010;
      15'b010_100001100010 : VALUE=19'b0000000_101000010010;
      15'b010_100001100011 : VALUE=19'b0000000_101000010010;
      15'b010_100001100100 : VALUE=19'b0000000_101000010010;
      15'b010_100001100101 : VALUE=19'b0000000_101000010010;
      15'b010_100001100110 : VALUE=19'b0000000_101000010010;
      15'b010_100001100111 : VALUE=19'b0000000_101000010010;
      15'b010_100001101000 : VALUE=19'b0000000_101000010001;
      15'b010_100001101001 : VALUE=19'b0000000_101000010001;
      15'b010_100001101010 : VALUE=19'b0000000_101000010001;
      15'b010_100001101011 : VALUE=19'b0000000_101000010001;
      15'b010_100001101100 : VALUE=19'b0000000_101000010001;
      15'b010_100001101101 : VALUE=19'b0000000_101000010001;
      15'b010_100001101110 : VALUE=19'b0000000_101000010001;
      15'b010_100001101111 : VALUE=19'b0000000_101000010001;
      15'b010_100001110000 : VALUE=19'b0000000_101000010000;
      15'b010_100001110001 : VALUE=19'b0000000_101000010000;
      15'b010_100001110010 : VALUE=19'b0000000_101000010000;
      15'b010_100001110011 : VALUE=19'b0000000_101000010000;
      15'b010_100001110100 : VALUE=19'b0000000_101000010000;
      15'b010_100001110101 : VALUE=19'b0000000_101000010000;
      15'b010_100001110110 : VALUE=19'b0000000_101000010000;
      15'b010_100001110111 : VALUE=19'b0000000_101000010000;
      15'b010_100001111000 : VALUE=19'b0000000_101000001111;
      15'b010_100001111001 : VALUE=19'b0000000_101000001111;
      15'b010_100001111010 : VALUE=19'b0000000_101000001111;
      15'b010_100001111011 : VALUE=19'b0000000_101000001111;
      15'b010_100001111100 : VALUE=19'b0000000_101000001111;
      15'b010_100001111101 : VALUE=19'b0000000_101000001111;
      15'b010_100001111110 : VALUE=19'b0000000_101000001111;
      15'b010_100001111111 : VALUE=19'b0000000_101000001111;
      15'b010_100010000000 : VALUE=19'b0000000_101000001110;
      15'b010_100010000001 : VALUE=19'b0000000_101000001110;
      15'b010_100010000010 : VALUE=19'b0000000_101000001110;
      15'b010_100010000011 : VALUE=19'b0000000_101000001110;
      15'b010_100010000100 : VALUE=19'b0000000_101000001110;
      15'b010_100010000101 : VALUE=19'b0000000_101000001110;
      15'b010_100010000110 : VALUE=19'b0000000_101000001110;
      15'b010_100010000111 : VALUE=19'b0000000_101000001110;
      15'b010_100010001000 : VALUE=19'b0000000_101000001110;
      15'b010_100010001001 : VALUE=19'b0000000_101000001101;
      15'b010_100010001010 : VALUE=19'b0000000_101000001101;
      15'b010_100010001011 : VALUE=19'b0000000_101000001101;
      15'b010_100010001100 : VALUE=19'b0000000_101000001101;
      15'b010_100010001101 : VALUE=19'b0000000_101000001101;
      15'b010_100010001110 : VALUE=19'b0000000_101000001101;
      15'b010_100010001111 : VALUE=19'b0000000_101000001101;
      15'b010_100010010000 : VALUE=19'b0000000_101000001101;
      15'b010_100010010001 : VALUE=19'b0000000_101000001100;
      15'b010_100010010010 : VALUE=19'b0000000_101000001100;
      15'b010_100010010011 : VALUE=19'b0000000_101000001100;
      15'b010_100010010100 : VALUE=19'b0000000_101000001100;
      15'b010_100010010101 : VALUE=19'b0000000_101000001100;
      15'b010_100010010110 : VALUE=19'b0000000_101000001100;
      15'b010_100010010111 : VALUE=19'b0000000_101000001100;
      15'b010_100010011000 : VALUE=19'b0000000_101000001100;
      15'b010_100010011001 : VALUE=19'b0000000_101000001011;
      15'b010_100010011010 : VALUE=19'b0000000_101000001011;
      15'b010_100010011011 : VALUE=19'b0000000_101000001011;
      15'b010_100010011100 : VALUE=19'b0000000_101000001011;
      15'b010_100010011101 : VALUE=19'b0000000_101000001011;
      15'b010_100010011110 : VALUE=19'b0000000_101000001011;
      15'b010_100010011111 : VALUE=19'b0000000_101000001011;
      15'b010_100010100000 : VALUE=19'b0000000_101000001011;
      15'b010_100010100001 : VALUE=19'b0000000_101000001010;
      15'b010_100010100010 : VALUE=19'b0000000_101000001010;
      15'b010_100010100011 : VALUE=19'b0000000_101000001010;
      15'b010_100010100100 : VALUE=19'b0000000_101000001010;
      15'b010_100010100101 : VALUE=19'b0000000_101000001010;
      15'b010_100010100110 : VALUE=19'b0000000_101000001010;
      15'b010_100010100111 : VALUE=19'b0000000_101000001010;
      15'b010_100010101000 : VALUE=19'b0000000_101000001010;
      15'b010_100010101001 : VALUE=19'b0000000_101000001001;
      15'b010_100010101010 : VALUE=19'b0000000_101000001001;
      15'b010_100010101011 : VALUE=19'b0000000_101000001001;
      15'b010_100010101100 : VALUE=19'b0000000_101000001001;
      15'b010_100010101101 : VALUE=19'b0000000_101000001001;
      15'b010_100010101110 : VALUE=19'b0000000_101000001001;
      15'b010_100010101111 : VALUE=19'b0000000_101000001001;
      15'b010_100010110000 : VALUE=19'b0000000_101000001001;
      15'b010_100010110001 : VALUE=19'b0000000_101000001000;
      15'b010_100010110010 : VALUE=19'b0000000_101000001000;
      15'b010_100010110011 : VALUE=19'b0000000_101000001000;
      15'b010_100010110100 : VALUE=19'b0000000_101000001000;
      15'b010_100010110101 : VALUE=19'b0000000_101000001000;
      15'b010_100010110110 : VALUE=19'b0000000_101000001000;
      15'b010_100010110111 : VALUE=19'b0000000_101000001000;
      15'b010_100010111000 : VALUE=19'b0000000_101000001000;
      15'b010_100010111001 : VALUE=19'b0000000_101000000111;
      15'b010_100010111010 : VALUE=19'b0000000_101000000111;
      15'b010_100010111011 : VALUE=19'b0000000_101000000111;
      15'b010_100010111100 : VALUE=19'b0000000_101000000111;
      15'b010_100010111101 : VALUE=19'b0000000_101000000111;
      15'b010_100010111110 : VALUE=19'b0000000_101000000111;
      15'b010_100010111111 : VALUE=19'b0000000_101000000111;
      15'b010_100011000000 : VALUE=19'b0000000_101000000111;
      15'b010_100011000001 : VALUE=19'b0000000_101000000110;
      15'b010_100011000010 : VALUE=19'b0000000_101000000110;
      15'b010_100011000011 : VALUE=19'b0000000_101000000110;
      15'b010_100011000100 : VALUE=19'b0000000_101000000110;
      15'b010_100011000101 : VALUE=19'b0000000_101000000110;
      15'b010_100011000110 : VALUE=19'b0000000_101000000110;
      15'b010_100011000111 : VALUE=19'b0000000_101000000110;
      15'b010_100011001000 : VALUE=19'b0000000_101000000110;
      15'b010_100011001001 : VALUE=19'b0000000_101000000101;
      15'b010_100011001010 : VALUE=19'b0000000_101000000101;
      15'b010_100011001011 : VALUE=19'b0000000_101000000101;
      15'b010_100011001100 : VALUE=19'b0000000_101000000101;
      15'b010_100011001101 : VALUE=19'b0000000_101000000101;
      15'b010_100011001110 : VALUE=19'b0000000_101000000101;
      15'b010_100011001111 : VALUE=19'b0000000_101000000101;
      15'b010_100011010000 : VALUE=19'b0000000_101000000101;
      15'b010_100011010001 : VALUE=19'b0000000_101000000100;
      15'b010_100011010010 : VALUE=19'b0000000_101000000100;
      15'b010_100011010011 : VALUE=19'b0000000_101000000100;
      15'b010_100011010100 : VALUE=19'b0000000_101000000100;
      15'b010_100011010101 : VALUE=19'b0000000_101000000100;
      15'b010_100011010110 : VALUE=19'b0000000_101000000100;
      15'b010_100011010111 : VALUE=19'b0000000_101000000100;
      15'b010_100011011000 : VALUE=19'b0000000_101000000100;
      15'b010_100011011001 : VALUE=19'b0000000_101000000100;
      15'b010_100011011010 : VALUE=19'b0000000_101000000011;
      15'b010_100011011011 : VALUE=19'b0000000_101000000011;
      15'b010_100011011100 : VALUE=19'b0000000_101000000011;
      15'b010_100011011101 : VALUE=19'b0000000_101000000011;
      15'b010_100011011110 : VALUE=19'b0000000_101000000011;
      15'b010_100011011111 : VALUE=19'b0000000_101000000011;
      15'b010_100011100000 : VALUE=19'b0000000_101000000011;
      15'b010_100011100001 : VALUE=19'b0000000_101000000011;
      15'b010_100011100010 : VALUE=19'b0000000_101000000010;
      15'b010_100011100011 : VALUE=19'b0000000_101000000010;
      15'b010_100011100100 : VALUE=19'b0000000_101000000010;
      15'b010_100011100101 : VALUE=19'b0000000_101000000010;
      15'b010_100011100110 : VALUE=19'b0000000_101000000010;
      15'b010_100011100111 : VALUE=19'b0000000_101000000010;
      15'b010_100011101000 : VALUE=19'b0000000_101000000010;
      15'b010_100011101001 : VALUE=19'b0000000_101000000010;
      15'b010_100011101010 : VALUE=19'b0000000_101000000001;
      15'b010_100011101011 : VALUE=19'b0000000_101000000001;
      15'b010_100011101100 : VALUE=19'b0000000_101000000001;
      15'b010_100011101101 : VALUE=19'b0000000_101000000001;
      15'b010_100011101110 : VALUE=19'b0000000_101000000001;
      15'b010_100011101111 : VALUE=19'b0000000_101000000001;
      15'b010_100011110000 : VALUE=19'b0000000_101000000001;
      15'b010_100011110001 : VALUE=19'b0000000_101000000001;
      15'b010_100011110010 : VALUE=19'b0000000_101000000000;
      15'b010_100011110011 : VALUE=19'b0000000_101000000000;
      15'b010_100011110100 : VALUE=19'b0000000_101000000000;
      15'b010_100011110101 : VALUE=19'b0000000_101000000000;
      15'b010_100011110110 : VALUE=19'b0000000_101000000000;
      15'b010_100011110111 : VALUE=19'b0000000_101000000000;
      15'b010_100011111000 : VALUE=19'b0000000_101000000000;
      15'b010_100011111001 : VALUE=19'b0000000_101000000000;
      15'b010_100011111010 : VALUE=19'b0000000_100111111111;
      15'b010_100011111011 : VALUE=19'b0000000_100111111111;
      15'b010_100011111100 : VALUE=19'b0000000_100111111111;
      15'b010_100011111101 : VALUE=19'b0000000_100111111111;
      15'b010_100011111110 : VALUE=19'b0000000_100111111111;
      15'b010_100011111111 : VALUE=19'b0000000_100111111111;
      15'b010_100100000000 : VALUE=19'b0000000_100111111111;
      15'b010_100100000001 : VALUE=19'b0000000_100111111111;
      15'b010_100100000010 : VALUE=19'b0000000_100111111111;
      15'b010_100100000011 : VALUE=19'b0000000_100111111110;
      15'b010_100100000100 : VALUE=19'b0000000_100111111110;
      15'b010_100100000101 : VALUE=19'b0000000_100111111110;
      15'b010_100100000110 : VALUE=19'b0000000_100111111110;
      15'b010_100100000111 : VALUE=19'b0000000_100111111110;
      15'b010_100100001000 : VALUE=19'b0000000_100111111110;
      15'b010_100100001001 : VALUE=19'b0000000_100111111110;
      15'b010_100100001010 : VALUE=19'b0000000_100111111110;
      15'b010_100100001011 : VALUE=19'b0000000_100111111101;
      15'b010_100100001100 : VALUE=19'b0000000_100111111101;
      15'b010_100100001101 : VALUE=19'b0000000_100111111101;
      15'b010_100100001110 : VALUE=19'b0000000_100111111101;
      15'b010_100100001111 : VALUE=19'b0000000_100111111101;
      15'b010_100100010000 : VALUE=19'b0000000_100111111101;
      15'b010_100100010001 : VALUE=19'b0000000_100111111101;
      15'b010_100100010010 : VALUE=19'b0000000_100111111101;
      15'b010_100100010011 : VALUE=19'b0000000_100111111100;
      15'b010_100100010100 : VALUE=19'b0000000_100111111100;
      15'b010_100100010101 : VALUE=19'b0000000_100111111100;
      15'b010_100100010110 : VALUE=19'b0000000_100111111100;
      15'b010_100100010111 : VALUE=19'b0000000_100111111100;
      15'b010_100100011000 : VALUE=19'b0000000_100111111100;
      15'b010_100100011001 : VALUE=19'b0000000_100111111100;
      15'b010_100100011010 : VALUE=19'b0000000_100111111100;
      15'b010_100100011011 : VALUE=19'b0000000_100111111011;
      15'b010_100100011100 : VALUE=19'b0000000_100111111011;
      15'b010_100100011101 : VALUE=19'b0000000_100111111011;
      15'b010_100100011110 : VALUE=19'b0000000_100111111011;
      15'b010_100100011111 : VALUE=19'b0000000_100111111011;
      15'b010_100100100000 : VALUE=19'b0000000_100111111011;
      15'b010_100100100001 : VALUE=19'b0000000_100111111011;
      15'b010_100100100010 : VALUE=19'b0000000_100111111011;
      15'b010_100100100011 : VALUE=19'b0000000_100111111010;
      15'b010_100100100100 : VALUE=19'b0000000_100111111010;
      15'b010_100100100101 : VALUE=19'b0000000_100111111010;
      15'b010_100100100110 : VALUE=19'b0000000_100111111010;
      15'b010_100100100111 : VALUE=19'b0000000_100111111010;
      15'b010_100100101000 : VALUE=19'b0000000_100111111010;
      15'b010_100100101001 : VALUE=19'b0000000_100111111010;
      15'b010_100100101010 : VALUE=19'b0000000_100111111010;
      15'b010_100100101011 : VALUE=19'b0000000_100111111010;
      15'b010_100100101100 : VALUE=19'b0000000_100111111001;
      15'b010_100100101101 : VALUE=19'b0000000_100111111001;
      15'b010_100100101110 : VALUE=19'b0000000_100111111001;
      15'b010_100100101111 : VALUE=19'b0000000_100111111001;
      15'b010_100100110000 : VALUE=19'b0000000_100111111001;
      15'b010_100100110001 : VALUE=19'b0000000_100111111001;
      15'b010_100100110010 : VALUE=19'b0000000_100111111001;
      15'b010_100100110011 : VALUE=19'b0000000_100111111001;
      15'b010_100100110100 : VALUE=19'b0000000_100111111000;
      15'b010_100100110101 : VALUE=19'b0000000_100111111000;
      15'b010_100100110110 : VALUE=19'b0000000_100111111000;
      15'b010_100100110111 : VALUE=19'b0000000_100111111000;
      15'b010_100100111000 : VALUE=19'b0000000_100111111000;
      15'b010_100100111001 : VALUE=19'b0000000_100111111000;
      15'b010_100100111010 : VALUE=19'b0000000_100111111000;
      15'b010_100100111011 : VALUE=19'b0000000_100111111000;
      15'b010_100100111100 : VALUE=19'b0000000_100111110111;
      15'b010_100100111101 : VALUE=19'b0000000_100111110111;
      15'b010_100100111110 : VALUE=19'b0000000_100111110111;
      15'b010_100100111111 : VALUE=19'b0000000_100111110111;
      15'b010_100101000000 : VALUE=19'b0000000_100111110111;
      15'b010_100101000001 : VALUE=19'b0000000_100111110111;
      15'b010_100101000010 : VALUE=19'b0000000_100111110111;
      15'b010_100101000011 : VALUE=19'b0000000_100111110111;
      15'b010_100101000100 : VALUE=19'b0000000_100111110111;
      15'b010_100101000101 : VALUE=19'b0000000_100111110110;
      15'b010_100101000110 : VALUE=19'b0000000_100111110110;
      15'b010_100101000111 : VALUE=19'b0000000_100111110110;
      15'b010_100101001000 : VALUE=19'b0000000_100111110110;
      15'b010_100101001001 : VALUE=19'b0000000_100111110110;
      15'b010_100101001010 : VALUE=19'b0000000_100111110110;
      15'b010_100101001011 : VALUE=19'b0000000_100111110110;
      15'b010_100101001100 : VALUE=19'b0000000_100111110110;
      15'b010_100101001101 : VALUE=19'b0000000_100111110101;
      15'b010_100101001110 : VALUE=19'b0000000_100111110101;
      15'b010_100101001111 : VALUE=19'b0000000_100111110101;
      15'b010_100101010000 : VALUE=19'b0000000_100111110101;
      15'b010_100101010001 : VALUE=19'b0000000_100111110101;
      15'b010_100101010010 : VALUE=19'b0000000_100111110101;
      15'b010_100101010011 : VALUE=19'b0000000_100111110101;
      15'b010_100101010100 : VALUE=19'b0000000_100111110101;
      15'b010_100101010101 : VALUE=19'b0000000_100111110100;
      15'b010_100101010110 : VALUE=19'b0000000_100111110100;
      15'b010_100101010111 : VALUE=19'b0000000_100111110100;
      15'b010_100101011000 : VALUE=19'b0000000_100111110100;
      15'b010_100101011001 : VALUE=19'b0000000_100111110100;
      15'b010_100101011010 : VALUE=19'b0000000_100111110100;
      15'b010_100101011011 : VALUE=19'b0000000_100111110100;
      15'b010_100101011100 : VALUE=19'b0000000_100111110100;
      15'b010_100101011101 : VALUE=19'b0000000_100111110011;
      15'b010_100101011110 : VALUE=19'b0000000_100111110011;
      15'b010_100101011111 : VALUE=19'b0000000_100111110011;
      15'b010_100101100000 : VALUE=19'b0000000_100111110011;
      15'b010_100101100001 : VALUE=19'b0000000_100111110011;
      15'b010_100101100010 : VALUE=19'b0000000_100111110011;
      15'b010_100101100011 : VALUE=19'b0000000_100111110011;
      15'b010_100101100100 : VALUE=19'b0000000_100111110011;
      15'b010_100101100101 : VALUE=19'b0000000_100111110011;
      15'b010_100101100110 : VALUE=19'b0000000_100111110010;
      15'b010_100101100111 : VALUE=19'b0000000_100111110010;
      15'b010_100101101000 : VALUE=19'b0000000_100111110010;
      15'b010_100101101001 : VALUE=19'b0000000_100111110010;
      15'b010_100101101010 : VALUE=19'b0000000_100111110010;
      15'b010_100101101011 : VALUE=19'b0000000_100111110010;
      15'b010_100101101100 : VALUE=19'b0000000_100111110010;
      15'b010_100101101101 : VALUE=19'b0000000_100111110010;
      15'b010_100101101110 : VALUE=19'b0000000_100111110001;
      15'b010_100101101111 : VALUE=19'b0000000_100111110001;
      15'b010_100101110000 : VALUE=19'b0000000_100111110001;
      15'b010_100101110001 : VALUE=19'b0000000_100111110001;
      15'b010_100101110010 : VALUE=19'b0000000_100111110001;
      15'b010_100101110011 : VALUE=19'b0000000_100111110001;
      15'b010_100101110100 : VALUE=19'b0000000_100111110001;
      15'b010_100101110101 : VALUE=19'b0000000_100111110001;
      15'b010_100101110110 : VALUE=19'b0000000_100111110000;
      15'b010_100101110111 : VALUE=19'b0000000_100111110000;
      15'b010_100101111000 : VALUE=19'b0000000_100111110000;
      15'b010_100101111001 : VALUE=19'b0000000_100111110000;
      15'b010_100101111010 : VALUE=19'b0000000_100111110000;
      15'b010_100101111011 : VALUE=19'b0000000_100111110000;
      15'b010_100101111100 : VALUE=19'b0000000_100111110000;
      15'b010_100101111101 : VALUE=19'b0000000_100111110000;
      15'b010_100101111110 : VALUE=19'b0000000_100111110000;
      15'b010_100101111111 : VALUE=19'b0000000_100111101111;
      15'b010_100110000000 : VALUE=19'b0000000_100111101111;
      15'b010_100110000001 : VALUE=19'b0000000_100111101111;
      15'b010_100110000010 : VALUE=19'b0000000_100111101111;
      15'b010_100110000011 : VALUE=19'b0000000_100111101111;
      15'b010_100110000100 : VALUE=19'b0000000_100111101111;
      15'b010_100110000101 : VALUE=19'b0000000_100111101111;
      15'b010_100110000110 : VALUE=19'b0000000_100111101111;
      15'b010_100110000111 : VALUE=19'b0000000_100111101110;
      15'b010_100110001000 : VALUE=19'b0000000_100111101110;
      15'b010_100110001001 : VALUE=19'b0000000_100111101110;
      15'b010_100110001010 : VALUE=19'b0000000_100111101110;
      15'b010_100110001011 : VALUE=19'b0000000_100111101110;
      15'b010_100110001100 : VALUE=19'b0000000_100111101110;
      15'b010_100110001101 : VALUE=19'b0000000_100111101110;
      15'b010_100110001110 : VALUE=19'b0000000_100111101110;
      15'b010_100110001111 : VALUE=19'b0000000_100111101101;
      15'b010_100110010000 : VALUE=19'b0000000_100111101101;
      15'b010_100110010001 : VALUE=19'b0000000_100111101101;
      15'b010_100110010010 : VALUE=19'b0000000_100111101101;
      15'b010_100110010011 : VALUE=19'b0000000_100111101101;
      15'b010_100110010100 : VALUE=19'b0000000_100111101101;
      15'b010_100110010101 : VALUE=19'b0000000_100111101101;
      15'b010_100110010110 : VALUE=19'b0000000_100111101101;
      15'b010_100110010111 : VALUE=19'b0000000_100111101101;
      15'b010_100110011000 : VALUE=19'b0000000_100111101100;
      15'b010_100110011001 : VALUE=19'b0000000_100111101100;
      15'b010_100110011010 : VALUE=19'b0000000_100111101100;
      15'b010_100110011011 : VALUE=19'b0000000_100111101100;
      15'b010_100110011100 : VALUE=19'b0000000_100111101100;
      15'b010_100110011101 : VALUE=19'b0000000_100111101100;
      15'b010_100110011110 : VALUE=19'b0000000_100111101100;
      15'b010_100110011111 : VALUE=19'b0000000_100111101100;
      15'b010_100110100000 : VALUE=19'b0000000_100111101011;
      15'b010_100110100001 : VALUE=19'b0000000_100111101011;
      15'b010_100110100010 : VALUE=19'b0000000_100111101011;
      15'b010_100110100011 : VALUE=19'b0000000_100111101011;
      15'b010_100110100100 : VALUE=19'b0000000_100111101011;
      15'b010_100110100101 : VALUE=19'b0000000_100111101011;
      15'b010_100110100110 : VALUE=19'b0000000_100111101011;
      15'b010_100110100111 : VALUE=19'b0000000_100111101011;
      15'b010_100110101000 : VALUE=19'b0000000_100111101011;
      15'b010_100110101001 : VALUE=19'b0000000_100111101010;
      15'b010_100110101010 : VALUE=19'b0000000_100111101010;
      15'b010_100110101011 : VALUE=19'b0000000_100111101010;
      15'b010_100110101100 : VALUE=19'b0000000_100111101010;
      15'b010_100110101101 : VALUE=19'b0000000_100111101010;
      15'b010_100110101110 : VALUE=19'b0000000_100111101010;
      15'b010_100110101111 : VALUE=19'b0000000_100111101010;
      15'b010_100110110000 : VALUE=19'b0000000_100111101010;
      15'b010_100110110001 : VALUE=19'b0000000_100111101001;
      15'b010_100110110010 : VALUE=19'b0000000_100111101001;
      15'b010_100110110011 : VALUE=19'b0000000_100111101001;
      15'b010_100110110100 : VALUE=19'b0000000_100111101001;
      15'b010_100110110101 : VALUE=19'b0000000_100111101001;
      15'b010_100110110110 : VALUE=19'b0000000_100111101001;
      15'b010_100110110111 : VALUE=19'b0000000_100111101001;
      15'b010_100110111000 : VALUE=19'b0000000_100111101001;
      15'b010_100110111001 : VALUE=19'b0000000_100111101000;
      15'b010_100110111010 : VALUE=19'b0000000_100111101000;
      15'b010_100110111011 : VALUE=19'b0000000_100111101000;
      15'b010_100110111100 : VALUE=19'b0000000_100111101000;
      15'b010_100110111101 : VALUE=19'b0000000_100111101000;
      15'b010_100110111110 : VALUE=19'b0000000_100111101000;
      15'b010_100110111111 : VALUE=19'b0000000_100111101000;
      15'b010_100111000000 : VALUE=19'b0000000_100111101000;
      15'b010_100111000001 : VALUE=19'b0000000_100111101000;
      15'b010_100111000010 : VALUE=19'b0000000_100111100111;
      15'b010_100111000011 : VALUE=19'b0000000_100111100111;
      15'b010_100111000100 : VALUE=19'b0000000_100111100111;
      15'b010_100111000101 : VALUE=19'b0000000_100111100111;
      15'b010_100111000110 : VALUE=19'b0000000_100111100111;
      15'b010_100111000111 : VALUE=19'b0000000_100111100111;
      15'b010_100111001000 : VALUE=19'b0000000_100111100111;
      15'b010_100111001001 : VALUE=19'b0000000_100111100111;
      15'b010_100111001010 : VALUE=19'b0000000_100111100110;
      15'b010_100111001011 : VALUE=19'b0000000_100111100110;
      15'b010_100111001100 : VALUE=19'b0000000_100111100110;
      15'b010_100111001101 : VALUE=19'b0000000_100111100110;
      15'b010_100111001110 : VALUE=19'b0000000_100111100110;
      15'b010_100111001111 : VALUE=19'b0000000_100111100110;
      15'b010_100111010000 : VALUE=19'b0000000_100111100110;
      15'b010_100111010001 : VALUE=19'b0000000_100111100110;
      15'b010_100111010010 : VALUE=19'b0000000_100111100110;
      15'b010_100111010011 : VALUE=19'b0000000_100111100101;
      15'b010_100111010100 : VALUE=19'b0000000_100111100101;
      15'b010_100111010101 : VALUE=19'b0000000_100111100101;
      15'b010_100111010110 : VALUE=19'b0000000_100111100101;
      15'b010_100111010111 : VALUE=19'b0000000_100111100101;
      15'b010_100111011000 : VALUE=19'b0000000_100111100101;
      15'b010_100111011001 : VALUE=19'b0000000_100111100101;
      15'b010_100111011010 : VALUE=19'b0000000_100111100101;
      15'b010_100111011011 : VALUE=19'b0000000_100111100100;
      15'b010_100111011100 : VALUE=19'b0000000_100111100100;
      15'b010_100111011101 : VALUE=19'b0000000_100111100100;
      15'b010_100111011110 : VALUE=19'b0000000_100111100100;
      15'b010_100111011111 : VALUE=19'b0000000_100111100100;
      15'b010_100111100000 : VALUE=19'b0000000_100111100100;
      15'b010_100111100001 : VALUE=19'b0000000_100111100100;
      15'b010_100111100010 : VALUE=19'b0000000_100111100100;
      15'b010_100111100011 : VALUE=19'b0000000_100111100100;
      15'b010_100111100100 : VALUE=19'b0000000_100111100011;
      15'b010_100111100101 : VALUE=19'b0000000_100111100011;
      15'b010_100111100110 : VALUE=19'b0000000_100111100011;
      15'b010_100111100111 : VALUE=19'b0000000_100111100011;
      15'b010_100111101000 : VALUE=19'b0000000_100111100011;
      15'b010_100111101001 : VALUE=19'b0000000_100111100011;
      15'b010_100111101010 : VALUE=19'b0000000_100111100011;
      15'b010_100111101011 : VALUE=19'b0000000_100111100011;
      15'b010_100111101100 : VALUE=19'b0000000_100111100010;
      15'b010_100111101101 : VALUE=19'b0000000_100111100010;
      15'b010_100111101110 : VALUE=19'b0000000_100111100010;
      15'b010_100111101111 : VALUE=19'b0000000_100111100010;
      15'b010_100111110000 : VALUE=19'b0000000_100111100010;
      15'b010_100111110001 : VALUE=19'b0000000_100111100010;
      15'b010_100111110010 : VALUE=19'b0000000_100111100010;
      15'b010_100111110011 : VALUE=19'b0000000_100111100010;
      15'b010_100111110100 : VALUE=19'b0000000_100111100010;
      15'b010_100111110101 : VALUE=19'b0000000_100111100001;
      15'b010_100111110110 : VALUE=19'b0000000_100111100001;
      15'b010_100111110111 : VALUE=19'b0000000_100111100001;
      15'b010_100111111000 : VALUE=19'b0000000_100111100001;
      15'b010_100111111001 : VALUE=19'b0000000_100111100001;
      15'b010_100111111010 : VALUE=19'b0000000_100111100001;
      15'b010_100111111011 : VALUE=19'b0000000_100111100001;
      15'b010_100111111100 : VALUE=19'b0000000_100111100001;
      15'b010_100111111101 : VALUE=19'b0000000_100111100000;
      15'b010_100111111110 : VALUE=19'b0000000_100111100000;
      15'b010_100111111111 : VALUE=19'b0000000_100111100000;
      15'b010_101000000000 : VALUE=19'b0000000_100111100000;
      15'b010_101000000001 : VALUE=19'b0000000_100111100000;
      15'b010_101000000010 : VALUE=19'b0000000_100111100000;
      15'b010_101000000011 : VALUE=19'b0000000_100111100000;
      15'b010_101000000100 : VALUE=19'b0000000_100111100000;
      15'b010_101000000101 : VALUE=19'b0000000_100111100000;
      15'b010_101000000110 : VALUE=19'b0000000_100111011111;
      15'b010_101000000111 : VALUE=19'b0000000_100111011111;
      15'b010_101000001000 : VALUE=19'b0000000_100111011111;
      15'b010_101000001001 : VALUE=19'b0000000_100111011111;
      15'b010_101000001010 : VALUE=19'b0000000_100111011111;
      15'b010_101000001011 : VALUE=19'b0000000_100111011111;
      15'b010_101000001100 : VALUE=19'b0000000_100111011111;
      15'b010_101000001101 : VALUE=19'b0000000_100111011111;
      15'b010_101000001110 : VALUE=19'b0000000_100111011110;
      15'b010_101000001111 : VALUE=19'b0000000_100111011110;
      15'b010_101000010000 : VALUE=19'b0000000_100111011110;
      15'b010_101000010001 : VALUE=19'b0000000_100111011110;
      15'b010_101000010010 : VALUE=19'b0000000_100111011110;
      15'b010_101000010011 : VALUE=19'b0000000_100111011110;
      15'b010_101000010100 : VALUE=19'b0000000_100111011110;
      15'b010_101000010101 : VALUE=19'b0000000_100111011110;
      15'b010_101000010110 : VALUE=19'b0000000_100111011110;
      15'b010_101000010111 : VALUE=19'b0000000_100111011101;
      15'b010_101000011000 : VALUE=19'b0000000_100111011101;
      15'b010_101000011001 : VALUE=19'b0000000_100111011101;
      15'b010_101000011010 : VALUE=19'b0000000_100111011101;
      15'b010_101000011011 : VALUE=19'b0000000_100111011101;
      15'b010_101000011100 : VALUE=19'b0000000_100111011101;
      15'b010_101000011101 : VALUE=19'b0000000_100111011101;
      15'b010_101000011110 : VALUE=19'b0000000_100111011101;
      15'b010_101000011111 : VALUE=19'b0000000_100111011100;
      15'b010_101000100000 : VALUE=19'b0000000_100111011100;
      15'b010_101000100001 : VALUE=19'b0000000_100111011100;
      15'b010_101000100010 : VALUE=19'b0000000_100111011100;
      15'b010_101000100011 : VALUE=19'b0000000_100111011100;
      15'b010_101000100100 : VALUE=19'b0000000_100111011100;
      15'b010_101000100101 : VALUE=19'b0000000_100111011100;
      15'b010_101000100110 : VALUE=19'b0000000_100111011100;
      15'b010_101000100111 : VALUE=19'b0000000_100111011100;
      15'b010_101000101000 : VALUE=19'b0000000_100111011011;
      15'b010_101000101001 : VALUE=19'b0000000_100111011011;
      15'b010_101000101010 : VALUE=19'b0000000_100111011011;
      15'b010_101000101011 : VALUE=19'b0000000_100111011011;
      15'b010_101000101100 : VALUE=19'b0000000_100111011011;
      15'b010_101000101101 : VALUE=19'b0000000_100111011011;
      15'b010_101000101110 : VALUE=19'b0000000_100111011011;
      15'b010_101000101111 : VALUE=19'b0000000_100111011011;
      15'b010_101000110000 : VALUE=19'b0000000_100111011010;
      15'b010_101000110001 : VALUE=19'b0000000_100111011010;
      15'b010_101000110010 : VALUE=19'b0000000_100111011010;
      15'b010_101000110011 : VALUE=19'b0000000_100111011010;
      15'b010_101000110100 : VALUE=19'b0000000_100111011010;
      15'b010_101000110101 : VALUE=19'b0000000_100111011010;
      15'b010_101000110110 : VALUE=19'b0000000_100111011010;
      15'b010_101000110111 : VALUE=19'b0000000_100111011010;
      15'b010_101000111000 : VALUE=19'b0000000_100111011010;
      15'b010_101000111001 : VALUE=19'b0000000_100111011001;
      15'b010_101000111010 : VALUE=19'b0000000_100111011001;
      15'b010_101000111011 : VALUE=19'b0000000_100111011001;
      15'b010_101000111100 : VALUE=19'b0000000_100111011001;
      15'b010_101000111101 : VALUE=19'b0000000_100111011001;
      15'b010_101000111110 : VALUE=19'b0000000_100111011001;
      15'b010_101000111111 : VALUE=19'b0000000_100111011001;
      15'b010_101001000000 : VALUE=19'b0000000_100111011001;
      15'b010_101001000001 : VALUE=19'b0000000_100111011000;
      15'b010_101001000010 : VALUE=19'b0000000_100111011000;
      15'b010_101001000011 : VALUE=19'b0000000_100111011000;
      15'b010_101001000100 : VALUE=19'b0000000_100111011000;
      15'b010_101001000101 : VALUE=19'b0000000_100111011000;
      15'b010_101001000110 : VALUE=19'b0000000_100111011000;
      15'b010_101001000111 : VALUE=19'b0000000_100111011000;
      15'b010_101001001000 : VALUE=19'b0000000_100111011000;
      15'b010_101001001001 : VALUE=19'b0000000_100111011000;
      15'b010_101001001010 : VALUE=19'b0000000_100111010111;
      15'b010_101001001011 : VALUE=19'b0000000_100111010111;
      15'b010_101001001100 : VALUE=19'b0000000_100111010111;
      15'b010_101001001101 : VALUE=19'b0000000_100111010111;
      15'b010_101001001110 : VALUE=19'b0000000_100111010111;
      15'b010_101001001111 : VALUE=19'b0000000_100111010111;
      15'b010_101001010000 : VALUE=19'b0000000_100111010111;
      15'b010_101001010001 : VALUE=19'b0000000_100111010111;
      15'b010_101001010010 : VALUE=19'b0000000_100111010111;
      15'b010_101001010011 : VALUE=19'b0000000_100111010110;
      15'b010_101001010100 : VALUE=19'b0000000_100111010110;
      15'b010_101001010101 : VALUE=19'b0000000_100111010110;
      15'b010_101001010110 : VALUE=19'b0000000_100111010110;
      15'b010_101001010111 : VALUE=19'b0000000_100111010110;
      15'b010_101001011000 : VALUE=19'b0000000_100111010110;
      15'b010_101001011001 : VALUE=19'b0000000_100111010110;
      15'b010_101001011010 : VALUE=19'b0000000_100111010110;
      15'b010_101001011011 : VALUE=19'b0000000_100111010101;
      15'b010_101001011100 : VALUE=19'b0000000_100111010101;
      15'b010_101001011101 : VALUE=19'b0000000_100111010101;
      15'b010_101001011110 : VALUE=19'b0000000_100111010101;
      15'b010_101001011111 : VALUE=19'b0000000_100111010101;
      15'b010_101001100000 : VALUE=19'b0000000_100111010101;
      15'b010_101001100001 : VALUE=19'b0000000_100111010101;
      15'b010_101001100010 : VALUE=19'b0000000_100111010101;
      15'b010_101001100011 : VALUE=19'b0000000_100111010101;
      15'b010_101001100100 : VALUE=19'b0000000_100111010100;
      15'b010_101001100101 : VALUE=19'b0000000_100111010100;
      15'b010_101001100110 : VALUE=19'b0000000_100111010100;
      15'b010_101001100111 : VALUE=19'b0000000_100111010100;
      15'b010_101001101000 : VALUE=19'b0000000_100111010100;
      15'b010_101001101001 : VALUE=19'b0000000_100111010100;
      15'b010_101001101010 : VALUE=19'b0000000_100111010100;
      15'b010_101001101011 : VALUE=19'b0000000_100111010100;
      15'b010_101001101100 : VALUE=19'b0000000_100111010100;
      15'b010_101001101101 : VALUE=19'b0000000_100111010011;
      15'b010_101001101110 : VALUE=19'b0000000_100111010011;
      15'b010_101001101111 : VALUE=19'b0000000_100111010011;
      15'b010_101001110000 : VALUE=19'b0000000_100111010011;
      15'b010_101001110001 : VALUE=19'b0000000_100111010011;
      15'b010_101001110010 : VALUE=19'b0000000_100111010011;
      15'b010_101001110011 : VALUE=19'b0000000_100111010011;
      15'b010_101001110100 : VALUE=19'b0000000_100111010011;
      15'b010_101001110101 : VALUE=19'b0000000_100111010010;
      15'b010_101001110110 : VALUE=19'b0000000_100111010010;
      15'b010_101001110111 : VALUE=19'b0000000_100111010010;
      15'b010_101001111000 : VALUE=19'b0000000_100111010010;
      15'b010_101001111001 : VALUE=19'b0000000_100111010010;
      15'b010_101001111010 : VALUE=19'b0000000_100111010010;
      15'b010_101001111011 : VALUE=19'b0000000_100111010010;
      15'b010_101001111100 : VALUE=19'b0000000_100111010010;
      15'b010_101001111101 : VALUE=19'b0000000_100111010010;
      15'b010_101001111110 : VALUE=19'b0000000_100111010001;
      15'b010_101001111111 : VALUE=19'b0000000_100111010001;
      15'b010_101010000000 : VALUE=19'b0000000_100111010001;
      15'b010_101010000001 : VALUE=19'b0000000_100111010001;
      15'b010_101010000010 : VALUE=19'b0000000_100111010001;
      15'b010_101010000011 : VALUE=19'b0000000_100111010001;
      15'b010_101010000100 : VALUE=19'b0000000_100111010001;
      15'b010_101010000101 : VALUE=19'b0000000_100111010001;
      15'b010_101010000110 : VALUE=19'b0000000_100111010000;
      15'b010_101010000111 : VALUE=19'b0000000_100111010000;
      15'b010_101010001000 : VALUE=19'b0000000_100111010000;
      15'b010_101010001001 : VALUE=19'b0000000_100111010000;
      15'b010_101010001010 : VALUE=19'b0000000_100111010000;
      15'b010_101010001011 : VALUE=19'b0000000_100111010000;
      15'b010_101010001100 : VALUE=19'b0000000_100111010000;
      15'b010_101010001101 : VALUE=19'b0000000_100111010000;
      15'b010_101010001110 : VALUE=19'b0000000_100111010000;
      15'b010_101010001111 : VALUE=19'b0000000_100111001111;
      15'b010_101010010000 : VALUE=19'b0000000_100111001111;
      15'b010_101010010001 : VALUE=19'b0000000_100111001111;
      15'b010_101010010010 : VALUE=19'b0000000_100111001111;
      15'b010_101010010011 : VALUE=19'b0000000_100111001111;
      15'b010_101010010100 : VALUE=19'b0000000_100111001111;
      15'b010_101010010101 : VALUE=19'b0000000_100111001111;
      15'b010_101010010110 : VALUE=19'b0000000_100111001111;
      15'b010_101010010111 : VALUE=19'b0000000_100111001111;
      15'b010_101010011000 : VALUE=19'b0000000_100111001110;
      15'b010_101010011001 : VALUE=19'b0000000_100111001110;
      15'b010_101010011010 : VALUE=19'b0000000_100111001110;
      15'b010_101010011011 : VALUE=19'b0000000_100111001110;
      15'b010_101010011100 : VALUE=19'b0000000_100111001110;
      15'b010_101010011101 : VALUE=19'b0000000_100111001110;
      15'b010_101010011110 : VALUE=19'b0000000_100111001110;
      15'b010_101010011111 : VALUE=19'b0000000_100111001110;
      15'b010_101010100000 : VALUE=19'b0000000_100111001110;
      15'b010_101010100001 : VALUE=19'b0000000_100111001101;
      15'b010_101010100010 : VALUE=19'b0000000_100111001101;
      15'b010_101010100011 : VALUE=19'b0000000_100111001101;
      15'b010_101010100100 : VALUE=19'b0000000_100111001101;
      15'b010_101010100101 : VALUE=19'b0000000_100111001101;
      15'b010_101010100110 : VALUE=19'b0000000_100111001101;
      15'b010_101010100111 : VALUE=19'b0000000_100111001101;
      15'b010_101010101000 : VALUE=19'b0000000_100111001101;
      15'b010_101010101001 : VALUE=19'b0000000_100111001100;
      15'b010_101010101010 : VALUE=19'b0000000_100111001100;
      15'b010_101010101011 : VALUE=19'b0000000_100111001100;
      15'b010_101010101100 : VALUE=19'b0000000_100111001100;
      15'b010_101010101101 : VALUE=19'b0000000_100111001100;
      15'b010_101010101110 : VALUE=19'b0000000_100111001100;
      15'b010_101010101111 : VALUE=19'b0000000_100111001100;
      15'b010_101010110000 : VALUE=19'b0000000_100111001100;
      15'b010_101010110001 : VALUE=19'b0000000_100111001100;
      15'b010_101010110010 : VALUE=19'b0000000_100111001011;
      15'b010_101010110011 : VALUE=19'b0000000_100111001011;
      15'b010_101010110100 : VALUE=19'b0000000_100111001011;
      15'b010_101010110101 : VALUE=19'b0000000_100111001011;
      15'b010_101010110110 : VALUE=19'b0000000_100111001011;
      15'b010_101010110111 : VALUE=19'b0000000_100111001011;
      15'b010_101010111000 : VALUE=19'b0000000_100111001011;
      15'b010_101010111001 : VALUE=19'b0000000_100111001011;
      15'b010_101010111010 : VALUE=19'b0000000_100111001011;
      15'b010_101010111011 : VALUE=19'b0000000_100111001010;
      15'b010_101010111100 : VALUE=19'b0000000_100111001010;
      15'b010_101010111101 : VALUE=19'b0000000_100111001010;
      15'b010_101010111110 : VALUE=19'b0000000_100111001010;
      15'b010_101010111111 : VALUE=19'b0000000_100111001010;
      15'b010_101011000000 : VALUE=19'b0000000_100111001010;
      15'b010_101011000001 : VALUE=19'b0000000_100111001010;
      15'b010_101011000010 : VALUE=19'b0000000_100111001010;
      15'b010_101011000011 : VALUE=19'b0000000_100111001001;
      15'b010_101011000100 : VALUE=19'b0000000_100111001001;
      15'b010_101011000101 : VALUE=19'b0000000_100111001001;
      15'b010_101011000110 : VALUE=19'b0000000_100111001001;
      15'b010_101011000111 : VALUE=19'b0000000_100111001001;
      15'b010_101011001000 : VALUE=19'b0000000_100111001001;
      15'b010_101011001001 : VALUE=19'b0000000_100111001001;
      15'b010_101011001010 : VALUE=19'b0000000_100111001001;
      15'b010_101011001011 : VALUE=19'b0000000_100111001001;
      15'b010_101011001100 : VALUE=19'b0000000_100111001000;
      15'b010_101011001101 : VALUE=19'b0000000_100111001000;
      15'b010_101011001110 : VALUE=19'b0000000_100111001000;
      15'b010_101011001111 : VALUE=19'b0000000_100111001000;
      15'b010_101011010000 : VALUE=19'b0000000_100111001000;
      15'b010_101011010001 : VALUE=19'b0000000_100111001000;
      15'b010_101011010010 : VALUE=19'b0000000_100111001000;
      15'b010_101011010011 : VALUE=19'b0000000_100111001000;
      15'b010_101011010100 : VALUE=19'b0000000_100111001000;
      15'b010_101011010101 : VALUE=19'b0000000_100111000111;
      15'b010_101011010110 : VALUE=19'b0000000_100111000111;
      15'b010_101011010111 : VALUE=19'b0000000_100111000111;
      15'b010_101011011000 : VALUE=19'b0000000_100111000111;
      15'b010_101011011001 : VALUE=19'b0000000_100111000111;
      15'b010_101011011010 : VALUE=19'b0000000_100111000111;
      15'b010_101011011011 : VALUE=19'b0000000_100111000111;
      15'b010_101011011100 : VALUE=19'b0000000_100111000111;
      15'b010_101011011101 : VALUE=19'b0000000_100111000111;
      15'b010_101011011110 : VALUE=19'b0000000_100111000110;
      15'b010_101011011111 : VALUE=19'b0000000_100111000110;
      15'b010_101011100000 : VALUE=19'b0000000_100111000110;
      15'b010_101011100001 : VALUE=19'b0000000_100111000110;
      15'b010_101011100010 : VALUE=19'b0000000_100111000110;
      15'b010_101011100011 : VALUE=19'b0000000_100111000110;
      15'b010_101011100100 : VALUE=19'b0000000_100111000110;
      15'b010_101011100101 : VALUE=19'b0000000_100111000110;
      15'b010_101011100110 : VALUE=19'b0000000_100111000101;
      15'b010_101011100111 : VALUE=19'b0000000_100111000101;
      15'b010_101011101000 : VALUE=19'b0000000_100111000101;
      15'b010_101011101001 : VALUE=19'b0000000_100111000101;
      15'b010_101011101010 : VALUE=19'b0000000_100111000101;
      15'b010_101011101011 : VALUE=19'b0000000_100111000101;
      15'b010_101011101100 : VALUE=19'b0000000_100111000101;
      15'b010_101011101101 : VALUE=19'b0000000_100111000101;
      15'b010_101011101110 : VALUE=19'b0000000_100111000101;
      15'b010_101011101111 : VALUE=19'b0000000_100111000100;
      15'b010_101011110000 : VALUE=19'b0000000_100111000100;
      15'b010_101011110001 : VALUE=19'b0000000_100111000100;
      15'b010_101011110010 : VALUE=19'b0000000_100111000100;
      15'b010_101011110011 : VALUE=19'b0000000_100111000100;
      15'b010_101011110100 : VALUE=19'b0000000_100111000100;
      15'b010_101011110101 : VALUE=19'b0000000_100111000100;
      15'b010_101011110110 : VALUE=19'b0000000_100111000100;
      15'b010_101011110111 : VALUE=19'b0000000_100111000100;
      15'b010_101011111000 : VALUE=19'b0000000_100111000011;
      15'b010_101011111001 : VALUE=19'b0000000_100111000011;
      15'b010_101011111010 : VALUE=19'b0000000_100111000011;
      15'b010_101011111011 : VALUE=19'b0000000_100111000011;
      15'b010_101011111100 : VALUE=19'b0000000_100111000011;
      15'b010_101011111101 : VALUE=19'b0000000_100111000011;
      15'b010_101011111110 : VALUE=19'b0000000_100111000011;
      15'b010_101011111111 : VALUE=19'b0000000_100111000011;
      15'b010_101100000000 : VALUE=19'b0000000_100111000011;
      15'b010_101100000001 : VALUE=19'b0000000_100111000010;
      15'b010_101100000010 : VALUE=19'b0000000_100111000010;
      15'b010_101100000011 : VALUE=19'b0000000_100111000010;
      15'b010_101100000100 : VALUE=19'b0000000_100111000010;
      15'b010_101100000101 : VALUE=19'b0000000_100111000010;
      15'b010_101100000110 : VALUE=19'b0000000_100111000010;
      15'b010_101100000111 : VALUE=19'b0000000_100111000010;
      15'b010_101100001000 : VALUE=19'b0000000_100111000010;
      15'b010_101100001001 : VALUE=19'b0000000_100111000010;
      15'b010_101100001010 : VALUE=19'b0000000_100111000001;
      15'b010_101100001011 : VALUE=19'b0000000_100111000001;
      15'b010_101100001100 : VALUE=19'b0000000_100111000001;
      15'b010_101100001101 : VALUE=19'b0000000_100111000001;
      15'b010_101100001110 : VALUE=19'b0000000_100111000001;
      15'b010_101100001111 : VALUE=19'b0000000_100111000001;
      15'b010_101100010000 : VALUE=19'b0000000_100111000001;
      15'b010_101100010001 : VALUE=19'b0000000_100111000001;
      15'b010_101100010010 : VALUE=19'b0000000_100111000000;
      15'b010_101100010011 : VALUE=19'b0000000_100111000000;
      15'b010_101100010100 : VALUE=19'b0000000_100111000000;
      15'b010_101100010101 : VALUE=19'b0000000_100111000000;
      15'b010_101100010110 : VALUE=19'b0000000_100111000000;
      15'b010_101100010111 : VALUE=19'b0000000_100111000000;
      15'b010_101100011000 : VALUE=19'b0000000_100111000000;
      15'b010_101100011001 : VALUE=19'b0000000_100111000000;
      15'b010_101100011010 : VALUE=19'b0000000_100111000000;
      15'b010_101100011011 : VALUE=19'b0000000_100110111111;
      15'b010_101100011100 : VALUE=19'b0000000_100110111111;
      15'b010_101100011101 : VALUE=19'b0000000_100110111111;
      15'b010_101100011110 : VALUE=19'b0000000_100110111111;
      15'b010_101100011111 : VALUE=19'b0000000_100110111111;
      15'b010_101100100000 : VALUE=19'b0000000_100110111111;
      15'b010_101100100001 : VALUE=19'b0000000_100110111111;
      15'b010_101100100010 : VALUE=19'b0000000_100110111111;
      15'b010_101100100011 : VALUE=19'b0000000_100110111111;
      15'b010_101100100100 : VALUE=19'b0000000_100110111110;
      15'b010_101100100101 : VALUE=19'b0000000_100110111110;
      15'b010_101100100110 : VALUE=19'b0000000_100110111110;
      15'b010_101100100111 : VALUE=19'b0000000_100110111110;
      15'b010_101100101000 : VALUE=19'b0000000_100110111110;
      15'b010_101100101001 : VALUE=19'b0000000_100110111110;
      15'b010_101100101010 : VALUE=19'b0000000_100110111110;
      15'b010_101100101011 : VALUE=19'b0000000_100110111110;
      15'b010_101100101100 : VALUE=19'b0000000_100110111110;
      15'b010_101100101101 : VALUE=19'b0000000_100110111101;
      15'b010_101100101110 : VALUE=19'b0000000_100110111101;
      15'b010_101100101111 : VALUE=19'b0000000_100110111101;
      15'b010_101100110000 : VALUE=19'b0000000_100110111101;
      15'b010_101100110001 : VALUE=19'b0000000_100110111101;
      15'b010_101100110010 : VALUE=19'b0000000_100110111101;
      15'b010_101100110011 : VALUE=19'b0000000_100110111101;
      15'b010_101100110100 : VALUE=19'b0000000_100110111101;
      15'b010_101100110101 : VALUE=19'b0000000_100110111101;
      15'b010_101100110110 : VALUE=19'b0000000_100110111100;
      15'b010_101100110111 : VALUE=19'b0000000_100110111100;
      15'b010_101100111000 : VALUE=19'b0000000_100110111100;
      15'b010_101100111001 : VALUE=19'b0000000_100110111100;
      15'b010_101100111010 : VALUE=19'b0000000_100110111100;
      15'b010_101100111011 : VALUE=19'b0000000_100110111100;
      15'b010_101100111100 : VALUE=19'b0000000_100110111100;
      15'b010_101100111101 : VALUE=19'b0000000_100110111100;
      15'b010_101100111110 : VALUE=19'b0000000_100110111100;
      15'b010_101100111111 : VALUE=19'b0000000_100110111011;
      15'b010_101101000000 : VALUE=19'b0000000_100110111011;
      15'b010_101101000001 : VALUE=19'b0000000_100110111011;
      15'b010_101101000010 : VALUE=19'b0000000_100110111011;
      15'b010_101101000011 : VALUE=19'b0000000_100110111011;
      15'b010_101101000100 : VALUE=19'b0000000_100110111011;
      15'b010_101101000101 : VALUE=19'b0000000_100110111011;
      15'b010_101101000110 : VALUE=19'b0000000_100110111011;
      15'b010_101101000111 : VALUE=19'b0000000_100110111011;
      15'b010_101101001000 : VALUE=19'b0000000_100110111010;
      15'b010_101101001001 : VALUE=19'b0000000_100110111010;
      15'b010_101101001010 : VALUE=19'b0000000_100110111010;
      15'b010_101101001011 : VALUE=19'b0000000_100110111010;
      15'b010_101101001100 : VALUE=19'b0000000_100110111010;
      15'b010_101101001101 : VALUE=19'b0000000_100110111010;
      15'b010_101101001110 : VALUE=19'b0000000_100110111010;
      15'b010_101101001111 : VALUE=19'b0000000_100110111010;
      15'b010_101101010000 : VALUE=19'b0000000_100110111010;
      15'b010_101101010001 : VALUE=19'b0000000_100110111001;
      15'b010_101101010010 : VALUE=19'b0000000_100110111001;
      15'b010_101101010011 : VALUE=19'b0000000_100110111001;
      15'b010_101101010100 : VALUE=19'b0000000_100110111001;
      15'b010_101101010101 : VALUE=19'b0000000_100110111001;
      15'b010_101101010110 : VALUE=19'b0000000_100110111001;
      15'b010_101101010111 : VALUE=19'b0000000_100110111001;
      15'b010_101101011000 : VALUE=19'b0000000_100110111001;
      15'b010_101101011001 : VALUE=19'b0000000_100110111000;
      15'b010_101101011010 : VALUE=19'b0000000_100110111000;
      15'b010_101101011011 : VALUE=19'b0000000_100110111000;
      15'b010_101101011100 : VALUE=19'b0000000_100110111000;
      15'b010_101101011101 : VALUE=19'b0000000_100110111000;
      15'b010_101101011110 : VALUE=19'b0000000_100110111000;
      15'b010_101101011111 : VALUE=19'b0000000_100110111000;
      15'b010_101101100000 : VALUE=19'b0000000_100110111000;
      15'b010_101101100001 : VALUE=19'b0000000_100110111000;
      15'b010_101101100010 : VALUE=19'b0000000_100110110111;
      15'b010_101101100011 : VALUE=19'b0000000_100110110111;
      15'b010_101101100100 : VALUE=19'b0000000_100110110111;
      15'b010_101101100101 : VALUE=19'b0000000_100110110111;
      15'b010_101101100110 : VALUE=19'b0000000_100110110111;
      15'b010_101101100111 : VALUE=19'b0000000_100110110111;
      15'b010_101101101000 : VALUE=19'b0000000_100110110111;
      15'b010_101101101001 : VALUE=19'b0000000_100110110111;
      15'b010_101101101010 : VALUE=19'b0000000_100110110111;
      15'b010_101101101011 : VALUE=19'b0000000_100110110110;
      15'b010_101101101100 : VALUE=19'b0000000_100110110110;
      15'b010_101101101101 : VALUE=19'b0000000_100110110110;
      15'b010_101101101110 : VALUE=19'b0000000_100110110110;
      15'b010_101101101111 : VALUE=19'b0000000_100110110110;
      15'b010_101101110000 : VALUE=19'b0000000_100110110110;
      15'b010_101101110001 : VALUE=19'b0000000_100110110110;
      15'b010_101101110010 : VALUE=19'b0000000_100110110110;
      15'b010_101101110011 : VALUE=19'b0000000_100110110110;
      15'b010_101101110100 : VALUE=19'b0000000_100110110101;
      15'b010_101101110101 : VALUE=19'b0000000_100110110101;
      15'b010_101101110110 : VALUE=19'b0000000_100110110101;
      15'b010_101101110111 : VALUE=19'b0000000_100110110101;
      15'b010_101101111000 : VALUE=19'b0000000_100110110101;
      15'b010_101101111001 : VALUE=19'b0000000_100110110101;
      15'b010_101101111010 : VALUE=19'b0000000_100110110101;
      15'b010_101101111011 : VALUE=19'b0000000_100110110101;
      15'b010_101101111100 : VALUE=19'b0000000_100110110101;
      15'b010_101101111101 : VALUE=19'b0000000_100110110100;
      15'b010_101101111110 : VALUE=19'b0000000_100110110100;
      15'b010_101101111111 : VALUE=19'b0000000_100110110100;
      15'b010_101110000000 : VALUE=19'b0000000_100110110100;
      15'b010_101110000001 : VALUE=19'b0000000_100110110100;
      15'b010_101110000010 : VALUE=19'b0000000_100110110100;
      15'b010_101110000011 : VALUE=19'b0000000_100110110100;
      15'b010_101110000100 : VALUE=19'b0000000_100110110100;
      15'b010_101110000101 : VALUE=19'b0000000_100110110100;
      15'b010_101110000110 : VALUE=19'b0000000_100110110011;
      15'b010_101110000111 : VALUE=19'b0000000_100110110011;
      15'b010_101110001000 : VALUE=19'b0000000_100110110011;
      15'b010_101110001001 : VALUE=19'b0000000_100110110011;
      15'b010_101110001010 : VALUE=19'b0000000_100110110011;
      15'b010_101110001011 : VALUE=19'b0000000_100110110011;
      15'b010_101110001100 : VALUE=19'b0000000_100110110011;
      15'b010_101110001101 : VALUE=19'b0000000_100110110011;
      15'b010_101110001110 : VALUE=19'b0000000_100110110011;
      15'b010_101110001111 : VALUE=19'b0000000_100110110010;
      15'b010_101110010000 : VALUE=19'b0000000_100110110010;
      15'b010_101110010001 : VALUE=19'b0000000_100110110010;
      15'b010_101110010010 : VALUE=19'b0000000_100110110010;
      15'b010_101110010011 : VALUE=19'b0000000_100110110010;
      15'b010_101110010100 : VALUE=19'b0000000_100110110010;
      15'b010_101110010101 : VALUE=19'b0000000_100110110010;
      15'b010_101110010110 : VALUE=19'b0000000_100110110010;
      15'b010_101110010111 : VALUE=19'b0000000_100110110010;
      15'b010_101110011000 : VALUE=19'b0000000_100110110001;
      15'b010_101110011001 : VALUE=19'b0000000_100110110001;
      15'b010_101110011010 : VALUE=19'b0000000_100110110001;
      15'b010_101110011011 : VALUE=19'b0000000_100110110001;
      15'b010_101110011100 : VALUE=19'b0000000_100110110001;
      15'b010_101110011101 : VALUE=19'b0000000_100110110001;
      15'b010_101110011110 : VALUE=19'b0000000_100110110001;
      15'b010_101110011111 : VALUE=19'b0000000_100110110001;
      15'b010_101110100000 : VALUE=19'b0000000_100110110001;
      15'b010_101110100001 : VALUE=19'b0000000_100110110000;
      15'b010_101110100010 : VALUE=19'b0000000_100110110000;
      15'b010_101110100011 : VALUE=19'b0000000_100110110000;
      15'b010_101110100100 : VALUE=19'b0000000_100110110000;
      15'b010_101110100101 : VALUE=19'b0000000_100110110000;
      15'b010_101110100110 : VALUE=19'b0000000_100110110000;
      15'b010_101110100111 : VALUE=19'b0000000_100110110000;
      15'b010_101110101000 : VALUE=19'b0000000_100110110000;
      15'b010_101110101001 : VALUE=19'b0000000_100110110000;
      15'b010_101110101010 : VALUE=19'b0000000_100110101111;
      15'b010_101110101011 : VALUE=19'b0000000_100110101111;
      15'b010_101110101100 : VALUE=19'b0000000_100110101111;
      15'b010_101110101101 : VALUE=19'b0000000_100110101111;
      15'b010_101110101110 : VALUE=19'b0000000_100110101111;
      15'b010_101110101111 : VALUE=19'b0000000_100110101111;
      15'b010_101110110000 : VALUE=19'b0000000_100110101111;
      15'b010_101110110001 : VALUE=19'b0000000_100110101111;
      15'b010_101110110010 : VALUE=19'b0000000_100110101111;
      15'b010_101110110011 : VALUE=19'b0000000_100110101110;
      15'b010_101110110100 : VALUE=19'b0000000_100110101110;
      15'b010_101110110101 : VALUE=19'b0000000_100110101110;
      15'b010_101110110110 : VALUE=19'b0000000_100110101110;
      15'b010_101110110111 : VALUE=19'b0000000_100110101110;
      15'b010_101110111000 : VALUE=19'b0000000_100110101110;
      15'b010_101110111001 : VALUE=19'b0000000_100110101110;
      15'b010_101110111010 : VALUE=19'b0000000_100110101110;
      15'b010_101110111011 : VALUE=19'b0000000_100110101110;
      15'b010_101110111100 : VALUE=19'b0000000_100110101101;
      15'b010_101110111101 : VALUE=19'b0000000_100110101101;
      15'b010_101110111110 : VALUE=19'b0000000_100110101101;
      15'b010_101110111111 : VALUE=19'b0000000_100110101101;
      15'b010_101111000000 : VALUE=19'b0000000_100110101101;
      15'b010_101111000001 : VALUE=19'b0000000_100110101101;
      15'b010_101111000010 : VALUE=19'b0000000_100110101101;
      15'b010_101111000011 : VALUE=19'b0000000_100110101101;
      15'b010_101111000100 : VALUE=19'b0000000_100110101101;
      15'b010_101111000101 : VALUE=19'b0000000_100110101100;
      15'b010_101111000110 : VALUE=19'b0000000_100110101100;
      15'b010_101111000111 : VALUE=19'b0000000_100110101100;
      15'b010_101111001000 : VALUE=19'b0000000_100110101100;
      15'b010_101111001001 : VALUE=19'b0000000_100110101100;
      15'b010_101111001010 : VALUE=19'b0000000_100110101100;
      15'b010_101111001011 : VALUE=19'b0000000_100110101100;
      15'b010_101111001100 : VALUE=19'b0000000_100110101100;
      15'b010_101111001101 : VALUE=19'b0000000_100110101100;
      15'b010_101111001110 : VALUE=19'b0000000_100110101011;
      15'b010_101111001111 : VALUE=19'b0000000_100110101011;
      15'b010_101111010000 : VALUE=19'b0000000_100110101011;
      15'b010_101111010001 : VALUE=19'b0000000_100110101011;
      15'b010_101111010010 : VALUE=19'b0000000_100110101011;
      15'b010_101111010011 : VALUE=19'b0000000_100110101011;
      15'b010_101111010100 : VALUE=19'b0000000_100110101011;
      15'b010_101111010101 : VALUE=19'b0000000_100110101011;
      15'b010_101111010110 : VALUE=19'b0000000_100110101011;
      15'b010_101111010111 : VALUE=19'b0000000_100110101010;
      15'b010_101111011000 : VALUE=19'b0000000_100110101010;
      15'b010_101111011001 : VALUE=19'b0000000_100110101010;
      15'b010_101111011010 : VALUE=19'b0000000_100110101010;
      15'b010_101111011011 : VALUE=19'b0000000_100110101010;
      15'b010_101111011100 : VALUE=19'b0000000_100110101010;
      15'b010_101111011101 : VALUE=19'b0000000_100110101010;
      15'b010_101111011110 : VALUE=19'b0000000_100110101010;
      15'b010_101111011111 : VALUE=19'b0000000_100110101010;
      15'b010_101111100000 : VALUE=19'b0000000_100110101001;
      15'b010_101111100001 : VALUE=19'b0000000_100110101001;
      15'b010_101111100010 : VALUE=19'b0000000_100110101001;
      15'b010_101111100011 : VALUE=19'b0000000_100110101001;
      15'b010_101111100100 : VALUE=19'b0000000_100110101001;
      15'b010_101111100101 : VALUE=19'b0000000_100110101001;
      15'b010_101111100110 : VALUE=19'b0000000_100110101001;
      15'b010_101111100111 : VALUE=19'b0000000_100110101001;
      15'b010_101111101000 : VALUE=19'b0000000_100110101001;
      15'b010_101111101001 : VALUE=19'b0000000_100110101001;
      15'b010_101111101010 : VALUE=19'b0000000_100110101000;
      15'b010_101111101011 : VALUE=19'b0000000_100110101000;
      15'b010_101111101100 : VALUE=19'b0000000_100110101000;
      15'b010_101111101101 : VALUE=19'b0000000_100110101000;
      15'b010_101111101110 : VALUE=19'b0000000_100110101000;
      15'b010_101111101111 : VALUE=19'b0000000_100110101000;
      15'b010_101111110000 : VALUE=19'b0000000_100110101000;
      15'b010_101111110001 : VALUE=19'b0000000_100110101000;
      15'b010_101111110010 : VALUE=19'b0000000_100110101000;
      15'b010_101111110011 : VALUE=19'b0000000_100110100111;
      15'b010_101111110100 : VALUE=19'b0000000_100110100111;
      15'b010_101111110101 : VALUE=19'b0000000_100110100111;
      15'b010_101111110110 : VALUE=19'b0000000_100110100111;
      15'b010_101111110111 : VALUE=19'b0000000_100110100111;
      15'b010_101111111000 : VALUE=19'b0000000_100110100111;
      15'b010_101111111001 : VALUE=19'b0000000_100110100111;
      15'b010_101111111010 : VALUE=19'b0000000_100110100111;
      15'b010_101111111011 : VALUE=19'b0000000_100110100111;
      15'b010_101111111100 : VALUE=19'b0000000_100110100110;
      15'b010_101111111101 : VALUE=19'b0000000_100110100110;
      15'b010_101111111110 : VALUE=19'b0000000_100110100110;
      15'b010_101111111111 : VALUE=19'b0000000_100110100110;
      15'b010_110000000000 : VALUE=19'b0000000_100110100110;
      15'b010_110000000001 : VALUE=19'b0000000_100110100110;
      15'b010_110000000010 : VALUE=19'b0000000_100110100110;
      15'b010_110000000011 : VALUE=19'b0000000_100110100110;
      15'b010_110000000100 : VALUE=19'b0000000_100110100110;
      15'b010_110000000101 : VALUE=19'b0000000_100110100101;
      15'b010_110000000110 : VALUE=19'b0000000_100110100101;
      15'b010_110000000111 : VALUE=19'b0000000_100110100101;
      15'b010_110000001000 : VALUE=19'b0000000_100110100101;
      15'b010_110000001001 : VALUE=19'b0000000_100110100101;
      15'b010_110000001010 : VALUE=19'b0000000_100110100101;
      15'b010_110000001011 : VALUE=19'b0000000_100110100101;
      15'b010_110000001100 : VALUE=19'b0000000_100110100101;
      15'b010_110000001101 : VALUE=19'b0000000_100110100101;
      15'b010_110000001110 : VALUE=19'b0000000_100110100100;
      15'b010_110000001111 : VALUE=19'b0000000_100110100100;
      15'b010_110000010000 : VALUE=19'b0000000_100110100100;
      15'b010_110000010001 : VALUE=19'b0000000_100110100100;
      15'b010_110000010010 : VALUE=19'b0000000_100110100100;
      15'b010_110000010011 : VALUE=19'b0000000_100110100100;
      15'b010_110000010100 : VALUE=19'b0000000_100110100100;
      15'b010_110000010101 : VALUE=19'b0000000_100110100100;
      15'b010_110000010110 : VALUE=19'b0000000_100110100100;
      15'b010_110000010111 : VALUE=19'b0000000_100110100011;
      15'b010_110000011000 : VALUE=19'b0000000_100110100011;
      15'b010_110000011001 : VALUE=19'b0000000_100110100011;
      15'b010_110000011010 : VALUE=19'b0000000_100110100011;
      15'b010_110000011011 : VALUE=19'b0000000_100110100011;
      15'b010_110000011100 : VALUE=19'b0000000_100110100011;
      15'b010_110000011101 : VALUE=19'b0000000_100110100011;
      15'b010_110000011110 : VALUE=19'b0000000_100110100011;
      15'b010_110000011111 : VALUE=19'b0000000_100110100011;
      15'b010_110000100000 : VALUE=19'b0000000_100110100010;
      15'b010_110000100001 : VALUE=19'b0000000_100110100010;
      15'b010_110000100010 : VALUE=19'b0000000_100110100010;
      15'b010_110000100011 : VALUE=19'b0000000_100110100010;
      15'b010_110000100100 : VALUE=19'b0000000_100110100010;
      15'b010_110000100101 : VALUE=19'b0000000_100110100010;
      15'b010_110000100110 : VALUE=19'b0000000_100110100010;
      15'b010_110000100111 : VALUE=19'b0000000_100110100010;
      15'b010_110000101000 : VALUE=19'b0000000_100110100010;
      15'b010_110000101001 : VALUE=19'b0000000_100110100001;
      15'b010_110000101010 : VALUE=19'b0000000_100110100001;
      15'b010_110000101011 : VALUE=19'b0000000_100110100001;
      15'b010_110000101100 : VALUE=19'b0000000_100110100001;
      15'b010_110000101101 : VALUE=19'b0000000_100110100001;
      15'b010_110000101110 : VALUE=19'b0000000_100110100001;
      15'b010_110000101111 : VALUE=19'b0000000_100110100001;
      15'b010_110000110000 : VALUE=19'b0000000_100110100001;
      15'b010_110000110001 : VALUE=19'b0000000_100110100001;
      15'b010_110000110010 : VALUE=19'b0000000_100110100001;
      15'b010_110000110011 : VALUE=19'b0000000_100110100000;
      15'b010_110000110100 : VALUE=19'b0000000_100110100000;
      15'b010_110000110101 : VALUE=19'b0000000_100110100000;
      15'b010_110000110110 : VALUE=19'b0000000_100110100000;
      15'b010_110000110111 : VALUE=19'b0000000_100110100000;
      15'b010_110000111000 : VALUE=19'b0000000_100110100000;
      15'b010_110000111001 : VALUE=19'b0000000_100110100000;
      15'b010_110000111010 : VALUE=19'b0000000_100110100000;
      15'b010_110000111011 : VALUE=19'b0000000_100110100000;
      15'b010_110000111100 : VALUE=19'b0000000_100110011111;
      15'b010_110000111101 : VALUE=19'b0000000_100110011111;
      15'b010_110000111110 : VALUE=19'b0000000_100110011111;
      15'b010_110000111111 : VALUE=19'b0000000_100110011111;
      15'b010_110001000000 : VALUE=19'b0000000_100110011111;
      15'b010_110001000001 : VALUE=19'b0000000_100110011111;
      15'b010_110001000010 : VALUE=19'b0000000_100110011111;
      15'b010_110001000011 : VALUE=19'b0000000_100110011111;
      15'b010_110001000100 : VALUE=19'b0000000_100110011111;
      15'b010_110001000101 : VALUE=19'b0000000_100110011110;
      15'b010_110001000110 : VALUE=19'b0000000_100110011110;
      15'b010_110001000111 : VALUE=19'b0000000_100110011110;
      15'b010_110001001000 : VALUE=19'b0000000_100110011110;
      15'b010_110001001001 : VALUE=19'b0000000_100110011110;
      15'b010_110001001010 : VALUE=19'b0000000_100110011110;
      15'b010_110001001011 : VALUE=19'b0000000_100110011110;
      15'b010_110001001100 : VALUE=19'b0000000_100110011110;
      15'b010_110001001101 : VALUE=19'b0000000_100110011110;
      15'b010_110001001110 : VALUE=19'b0000000_100110011101;
      15'b010_110001001111 : VALUE=19'b0000000_100110011101;
      15'b010_110001010000 : VALUE=19'b0000000_100110011101;
      15'b010_110001010001 : VALUE=19'b0000000_100110011101;
      15'b010_110001010010 : VALUE=19'b0000000_100110011101;
      15'b010_110001010011 : VALUE=19'b0000000_100110011101;
      15'b010_110001010100 : VALUE=19'b0000000_100110011101;
      15'b010_110001010101 : VALUE=19'b0000000_100110011101;
      15'b010_110001010110 : VALUE=19'b0000000_100110011101;
      15'b010_110001010111 : VALUE=19'b0000000_100110011100;
      15'b010_110001011000 : VALUE=19'b0000000_100110011100;
      15'b010_110001011001 : VALUE=19'b0000000_100110011100;
      15'b010_110001011010 : VALUE=19'b0000000_100110011100;
      15'b010_110001011011 : VALUE=19'b0000000_100110011100;
      15'b010_110001011100 : VALUE=19'b0000000_100110011100;
      15'b010_110001011101 : VALUE=19'b0000000_100110011100;
      15'b010_110001011110 : VALUE=19'b0000000_100110011100;
      15'b010_110001011111 : VALUE=19'b0000000_100110011100;
      15'b010_110001100000 : VALUE=19'b0000000_100110011100;
      15'b010_110001100001 : VALUE=19'b0000000_100110011011;
      15'b010_110001100010 : VALUE=19'b0000000_100110011011;
      15'b010_110001100011 : VALUE=19'b0000000_100110011011;
      15'b010_110001100100 : VALUE=19'b0000000_100110011011;
      15'b010_110001100101 : VALUE=19'b0000000_100110011011;
      15'b010_110001100110 : VALUE=19'b0000000_100110011011;
      15'b010_110001100111 : VALUE=19'b0000000_100110011011;
      15'b010_110001101000 : VALUE=19'b0000000_100110011011;
      15'b010_110001101001 : VALUE=19'b0000000_100110011011;
      15'b010_110001101010 : VALUE=19'b0000000_100110011010;
      15'b010_110001101011 : VALUE=19'b0000000_100110011010;
      15'b010_110001101100 : VALUE=19'b0000000_100110011010;
      15'b010_110001101101 : VALUE=19'b0000000_100110011010;
      15'b010_110001101110 : VALUE=19'b0000000_100110011010;
      15'b010_110001101111 : VALUE=19'b0000000_100110011010;
      15'b010_110001110000 : VALUE=19'b0000000_100110011010;
      15'b010_110001110001 : VALUE=19'b0000000_100110011010;
      15'b010_110001110010 : VALUE=19'b0000000_100110011010;
      15'b010_110001110011 : VALUE=19'b0000000_100110011001;
      15'b010_110001110100 : VALUE=19'b0000000_100110011001;
      15'b010_110001110101 : VALUE=19'b0000000_100110011001;
      15'b010_110001110110 : VALUE=19'b0000000_100110011001;
      15'b010_110001110111 : VALUE=19'b0000000_100110011001;
      15'b010_110001111000 : VALUE=19'b0000000_100110011001;
      15'b010_110001111001 : VALUE=19'b0000000_100110011001;
      15'b010_110001111010 : VALUE=19'b0000000_100110011001;
      15'b010_110001111011 : VALUE=19'b0000000_100110011001;
      15'b010_110001111100 : VALUE=19'b0000000_100110011000;
      15'b010_110001111101 : VALUE=19'b0000000_100110011000;
      15'b010_110001111110 : VALUE=19'b0000000_100110011000;
      15'b010_110001111111 : VALUE=19'b0000000_100110011000;
      15'b010_110010000000 : VALUE=19'b0000000_100110011000;
      15'b010_110010000001 : VALUE=19'b0000000_100110011000;
      15'b010_110010000010 : VALUE=19'b0000000_100110011000;
      15'b010_110010000011 : VALUE=19'b0000000_100110011000;
      15'b010_110010000100 : VALUE=19'b0000000_100110011000;
      15'b010_110010000101 : VALUE=19'b0000000_100110011000;
      15'b010_110010000110 : VALUE=19'b0000000_100110010111;
      15'b010_110010000111 : VALUE=19'b0000000_100110010111;
      15'b010_110010001000 : VALUE=19'b0000000_100110010111;
      15'b010_110010001001 : VALUE=19'b0000000_100110010111;
      15'b010_110010001010 : VALUE=19'b0000000_100110010111;
      15'b010_110010001011 : VALUE=19'b0000000_100110010111;
      15'b010_110010001100 : VALUE=19'b0000000_100110010111;
      15'b010_110010001101 : VALUE=19'b0000000_100110010111;
      15'b010_110010001110 : VALUE=19'b0000000_100110010111;
      15'b010_110010001111 : VALUE=19'b0000000_100110010110;
      15'b010_110010010000 : VALUE=19'b0000000_100110010110;
      15'b010_110010010001 : VALUE=19'b0000000_100110010110;
      15'b010_110010010010 : VALUE=19'b0000000_100110010110;
      15'b010_110010010011 : VALUE=19'b0000000_100110010110;
      15'b010_110010010100 : VALUE=19'b0000000_100110010110;
      15'b010_110010010101 : VALUE=19'b0000000_100110010110;
      15'b010_110010010110 : VALUE=19'b0000000_100110010110;
      15'b010_110010010111 : VALUE=19'b0000000_100110010110;
      15'b010_110010011000 : VALUE=19'b0000000_100110010101;
      15'b010_110010011001 : VALUE=19'b0000000_100110010101;
      15'b010_110010011010 : VALUE=19'b0000000_100110010101;
      15'b010_110010011011 : VALUE=19'b0000000_100110010101;
      15'b010_110010011100 : VALUE=19'b0000000_100110010101;
      15'b010_110010011101 : VALUE=19'b0000000_100110010101;
      15'b010_110010011110 : VALUE=19'b0000000_100110010101;
      15'b010_110010011111 : VALUE=19'b0000000_100110010101;
      15'b010_110010100000 : VALUE=19'b0000000_100110010101;
      15'b010_110010100001 : VALUE=19'b0000000_100110010101;
      15'b010_110010100010 : VALUE=19'b0000000_100110010100;
      15'b010_110010100011 : VALUE=19'b0000000_100110010100;
      15'b010_110010100100 : VALUE=19'b0000000_100110010100;
      15'b010_110010100101 : VALUE=19'b0000000_100110010100;
      15'b010_110010100110 : VALUE=19'b0000000_100110010100;
      15'b010_110010100111 : VALUE=19'b0000000_100110010100;
      15'b010_110010101000 : VALUE=19'b0000000_100110010100;
      15'b010_110010101001 : VALUE=19'b0000000_100110010100;
      15'b010_110010101010 : VALUE=19'b0000000_100110010100;
      15'b010_110010101011 : VALUE=19'b0000000_100110010011;
      15'b010_110010101100 : VALUE=19'b0000000_100110010011;
      15'b010_110010101101 : VALUE=19'b0000000_100110010011;
      15'b010_110010101110 : VALUE=19'b0000000_100110010011;
      15'b010_110010101111 : VALUE=19'b0000000_100110010011;
      15'b010_110010110000 : VALUE=19'b0000000_100110010011;
      15'b010_110010110001 : VALUE=19'b0000000_100110010011;
      15'b010_110010110010 : VALUE=19'b0000000_100110010011;
      15'b010_110010110011 : VALUE=19'b0000000_100110010011;
      15'b010_110010110100 : VALUE=19'b0000000_100110010010;
      15'b010_110010110101 : VALUE=19'b0000000_100110010010;
      15'b010_110010110110 : VALUE=19'b0000000_100110010010;
      15'b010_110010110111 : VALUE=19'b0000000_100110010010;
      15'b010_110010111000 : VALUE=19'b0000000_100110010010;
      15'b010_110010111001 : VALUE=19'b0000000_100110010010;
      15'b010_110010111010 : VALUE=19'b0000000_100110010010;
      15'b010_110010111011 : VALUE=19'b0000000_100110010010;
      15'b010_110010111100 : VALUE=19'b0000000_100110010010;
      15'b010_110010111101 : VALUE=19'b0000000_100110010010;
      15'b010_110010111110 : VALUE=19'b0000000_100110010001;
      15'b010_110010111111 : VALUE=19'b0000000_100110010001;
      15'b010_110011000000 : VALUE=19'b0000000_100110010001;
      15'b010_110011000001 : VALUE=19'b0000000_100110010001;
      15'b010_110011000010 : VALUE=19'b0000000_100110010001;
      15'b010_110011000011 : VALUE=19'b0000000_100110010001;
      15'b010_110011000100 : VALUE=19'b0000000_100110010001;
      15'b010_110011000101 : VALUE=19'b0000000_100110010001;
      15'b010_110011000110 : VALUE=19'b0000000_100110010001;
      15'b010_110011000111 : VALUE=19'b0000000_100110010000;
      15'b010_110011001000 : VALUE=19'b0000000_100110010000;
      15'b010_110011001001 : VALUE=19'b0000000_100110010000;
      15'b010_110011001010 : VALUE=19'b0000000_100110010000;
      15'b010_110011001011 : VALUE=19'b0000000_100110010000;
      15'b010_110011001100 : VALUE=19'b0000000_100110010000;
      15'b010_110011001101 : VALUE=19'b0000000_100110010000;
      15'b010_110011001110 : VALUE=19'b0000000_100110010000;
      15'b010_110011001111 : VALUE=19'b0000000_100110010000;
      15'b010_110011010000 : VALUE=19'b0000000_100110001111;
      15'b010_110011010001 : VALUE=19'b0000000_100110001111;
      15'b010_110011010010 : VALUE=19'b0000000_100110001111;
      15'b010_110011010011 : VALUE=19'b0000000_100110001111;
      15'b010_110011010100 : VALUE=19'b0000000_100110001111;
      15'b010_110011010101 : VALUE=19'b0000000_100110001111;
      15'b010_110011010110 : VALUE=19'b0000000_100110001111;
      15'b010_110011010111 : VALUE=19'b0000000_100110001111;
      15'b010_110011011000 : VALUE=19'b0000000_100110001111;
      15'b010_110011011001 : VALUE=19'b0000000_100110001111;
      15'b010_110011011010 : VALUE=19'b0000000_100110001110;
      15'b010_110011011011 : VALUE=19'b0000000_100110001110;
      15'b010_110011011100 : VALUE=19'b0000000_100110001110;
      15'b010_110011011101 : VALUE=19'b0000000_100110001110;
      15'b010_110011011110 : VALUE=19'b0000000_100110001110;
      15'b010_110011011111 : VALUE=19'b0000000_100110001110;
      15'b010_110011100000 : VALUE=19'b0000000_100110001110;
      15'b010_110011100001 : VALUE=19'b0000000_100110001110;
      15'b010_110011100010 : VALUE=19'b0000000_100110001110;
      15'b010_110011100011 : VALUE=19'b0000000_100110001101;
      15'b010_110011100100 : VALUE=19'b0000000_100110001101;
      15'b010_110011100101 : VALUE=19'b0000000_100110001101;
      15'b010_110011100110 : VALUE=19'b0000000_100110001101;
      15'b010_110011100111 : VALUE=19'b0000000_100110001101;
      15'b010_110011101000 : VALUE=19'b0000000_100110001101;
      15'b010_110011101001 : VALUE=19'b0000000_100110001101;
      15'b010_110011101010 : VALUE=19'b0000000_100110001101;
      15'b010_110011101011 : VALUE=19'b0000000_100110001101;
      15'b010_110011101100 : VALUE=19'b0000000_100110001101;
      15'b010_110011101101 : VALUE=19'b0000000_100110001100;
      15'b010_110011101110 : VALUE=19'b0000000_100110001100;
      15'b010_110011101111 : VALUE=19'b0000000_100110001100;
      15'b010_110011110000 : VALUE=19'b0000000_100110001100;
      15'b010_110011110001 : VALUE=19'b0000000_100110001100;
      15'b010_110011110010 : VALUE=19'b0000000_100110001100;
      15'b010_110011110011 : VALUE=19'b0000000_100110001100;
      15'b010_110011110100 : VALUE=19'b0000000_100110001100;
      15'b010_110011110101 : VALUE=19'b0000000_100110001100;
      15'b010_110011110110 : VALUE=19'b0000000_100110001011;
      15'b010_110011110111 : VALUE=19'b0000000_100110001011;
      15'b010_110011111000 : VALUE=19'b0000000_100110001011;
      15'b010_110011111001 : VALUE=19'b0000000_100110001011;
      15'b010_110011111010 : VALUE=19'b0000000_100110001011;
      15'b010_110011111011 : VALUE=19'b0000000_100110001011;
      15'b010_110011111100 : VALUE=19'b0000000_100110001011;
      15'b010_110011111101 : VALUE=19'b0000000_100110001011;
      15'b010_110011111110 : VALUE=19'b0000000_100110001011;
      15'b010_110011111111 : VALUE=19'b0000000_100110001010;
      15'b010_110100000000 : VALUE=19'b0000000_100110001010;
      15'b010_110100000001 : VALUE=19'b0000000_100110001010;
      15'b010_110100000010 : VALUE=19'b0000000_100110001010;
      15'b010_110100000011 : VALUE=19'b0000000_100110001010;
      15'b010_110100000100 : VALUE=19'b0000000_100110001010;
      15'b010_110100000101 : VALUE=19'b0000000_100110001010;
      15'b010_110100000110 : VALUE=19'b0000000_100110001010;
      15'b010_110100000111 : VALUE=19'b0000000_100110001010;
      15'b010_110100001000 : VALUE=19'b0000000_100110001010;
      15'b010_110100001001 : VALUE=19'b0000000_100110001001;
      15'b010_110100001010 : VALUE=19'b0000000_100110001001;
      15'b010_110100001011 : VALUE=19'b0000000_100110001001;
      15'b010_110100001100 : VALUE=19'b0000000_100110001001;
      15'b010_110100001101 : VALUE=19'b0000000_100110001001;
      15'b010_110100001110 : VALUE=19'b0000000_100110001001;
      15'b010_110100001111 : VALUE=19'b0000000_100110001001;
      15'b010_110100010000 : VALUE=19'b0000000_100110001001;
      15'b010_110100010001 : VALUE=19'b0000000_100110001001;
      15'b010_110100010010 : VALUE=19'b0000000_100110001000;
      15'b010_110100010011 : VALUE=19'b0000000_100110001000;
      15'b010_110100010100 : VALUE=19'b0000000_100110001000;
      15'b010_110100010101 : VALUE=19'b0000000_100110001000;
      15'b010_110100010110 : VALUE=19'b0000000_100110001000;
      15'b010_110100010111 : VALUE=19'b0000000_100110001000;
      15'b010_110100011000 : VALUE=19'b0000000_100110001000;
      15'b010_110100011001 : VALUE=19'b0000000_100110001000;
      15'b010_110100011010 : VALUE=19'b0000000_100110001000;
      15'b010_110100011011 : VALUE=19'b0000000_100110001000;
      15'b010_110100011100 : VALUE=19'b0000000_100110000111;
      15'b010_110100011101 : VALUE=19'b0000000_100110000111;
      15'b010_110100011110 : VALUE=19'b0000000_100110000111;
      15'b010_110100011111 : VALUE=19'b0000000_100110000111;
      15'b010_110100100000 : VALUE=19'b0000000_100110000111;
      15'b010_110100100001 : VALUE=19'b0000000_100110000111;
      15'b010_110100100010 : VALUE=19'b0000000_100110000111;
      15'b010_110100100011 : VALUE=19'b0000000_100110000111;
      15'b010_110100100100 : VALUE=19'b0000000_100110000111;
      15'b010_110100100101 : VALUE=19'b0000000_100110000110;
      15'b010_110100100110 : VALUE=19'b0000000_100110000110;
      15'b010_110100100111 : VALUE=19'b0000000_100110000110;
      15'b010_110100101000 : VALUE=19'b0000000_100110000110;
      15'b010_110100101001 : VALUE=19'b0000000_100110000110;
      15'b010_110100101010 : VALUE=19'b0000000_100110000110;
      15'b010_110100101011 : VALUE=19'b0000000_100110000110;
      15'b010_110100101100 : VALUE=19'b0000000_100110000110;
      15'b010_110100101101 : VALUE=19'b0000000_100110000110;
      15'b010_110100101110 : VALUE=19'b0000000_100110000110;
      15'b010_110100101111 : VALUE=19'b0000000_100110000101;
      15'b010_110100110000 : VALUE=19'b0000000_100110000101;
      15'b010_110100110001 : VALUE=19'b0000000_100110000101;
      15'b010_110100110010 : VALUE=19'b0000000_100110000101;
      15'b010_110100110011 : VALUE=19'b0000000_100110000101;
      15'b010_110100110100 : VALUE=19'b0000000_100110000101;
      15'b010_110100110101 : VALUE=19'b0000000_100110000101;
      15'b010_110100110110 : VALUE=19'b0000000_100110000101;
      15'b010_110100110111 : VALUE=19'b0000000_100110000101;
      15'b010_110100111000 : VALUE=19'b0000000_100110000100;
      15'b010_110100111001 : VALUE=19'b0000000_100110000100;
      15'b010_110100111010 : VALUE=19'b0000000_100110000100;
      15'b010_110100111011 : VALUE=19'b0000000_100110000100;
      15'b010_110100111100 : VALUE=19'b0000000_100110000100;
      15'b010_110100111101 : VALUE=19'b0000000_100110000100;
      15'b010_110100111110 : VALUE=19'b0000000_100110000100;
      15'b010_110100111111 : VALUE=19'b0000000_100110000100;
      15'b010_110101000000 : VALUE=19'b0000000_100110000100;
      15'b010_110101000001 : VALUE=19'b0000000_100110000100;
      15'b010_110101000010 : VALUE=19'b0000000_100110000011;
      15'b010_110101000011 : VALUE=19'b0000000_100110000011;
      15'b010_110101000100 : VALUE=19'b0000000_100110000011;
      15'b010_110101000101 : VALUE=19'b0000000_100110000011;
      15'b010_110101000110 : VALUE=19'b0000000_100110000011;
      15'b010_110101000111 : VALUE=19'b0000000_100110000011;
      15'b010_110101001000 : VALUE=19'b0000000_100110000011;
      15'b010_110101001001 : VALUE=19'b0000000_100110000011;
      15'b010_110101001010 : VALUE=19'b0000000_100110000011;
      15'b010_110101001011 : VALUE=19'b0000000_100110000010;
      15'b010_110101001100 : VALUE=19'b0000000_100110000010;
      15'b010_110101001101 : VALUE=19'b0000000_100110000010;
      15'b010_110101001110 : VALUE=19'b0000000_100110000010;
      15'b010_110101001111 : VALUE=19'b0000000_100110000010;
      15'b010_110101010000 : VALUE=19'b0000000_100110000010;
      15'b010_110101010001 : VALUE=19'b0000000_100110000010;
      15'b010_110101010010 : VALUE=19'b0000000_100110000010;
      15'b010_110101010011 : VALUE=19'b0000000_100110000010;
      15'b010_110101010100 : VALUE=19'b0000000_100110000010;
      15'b010_110101010101 : VALUE=19'b0000000_100110000001;
      15'b010_110101010110 : VALUE=19'b0000000_100110000001;
      15'b010_110101010111 : VALUE=19'b0000000_100110000001;
      15'b010_110101011000 : VALUE=19'b0000000_100110000001;
      15'b010_110101011001 : VALUE=19'b0000000_100110000001;
      15'b010_110101011010 : VALUE=19'b0000000_100110000001;
      15'b010_110101011011 : VALUE=19'b0000000_100110000001;
      15'b010_110101011100 : VALUE=19'b0000000_100110000001;
      15'b010_110101011101 : VALUE=19'b0000000_100110000001;
      15'b010_110101011110 : VALUE=19'b0000000_100110000000;
      15'b010_110101011111 : VALUE=19'b0000000_100110000000;
      15'b010_110101100000 : VALUE=19'b0000000_100110000000;
      15'b010_110101100001 : VALUE=19'b0000000_100110000000;
      15'b010_110101100010 : VALUE=19'b0000000_100110000000;
      15'b010_110101100011 : VALUE=19'b0000000_100110000000;
      15'b010_110101100100 : VALUE=19'b0000000_100110000000;
      15'b010_110101100101 : VALUE=19'b0000000_100110000000;
      15'b010_110101100110 : VALUE=19'b0000000_100110000000;
      15'b010_110101100111 : VALUE=19'b0000000_100110000000;
      15'b010_110101101000 : VALUE=19'b0000000_100101111111;
      15'b010_110101101001 : VALUE=19'b0000000_100101111111;
      15'b010_110101101010 : VALUE=19'b0000000_100101111111;
      15'b010_110101101011 : VALUE=19'b0000000_100101111111;
      15'b010_110101101100 : VALUE=19'b0000000_100101111111;
      15'b010_110101101101 : VALUE=19'b0000000_100101111111;
      15'b010_110101101110 : VALUE=19'b0000000_100101111111;
      15'b010_110101101111 : VALUE=19'b0000000_100101111111;
      15'b010_110101110000 : VALUE=19'b0000000_100101111111;
      15'b010_110101110001 : VALUE=19'b0000000_100101111110;
      15'b010_110101110010 : VALUE=19'b0000000_100101111110;
      15'b010_110101110011 : VALUE=19'b0000000_100101111110;
      15'b010_110101110100 : VALUE=19'b0000000_100101111110;
      15'b010_110101110101 : VALUE=19'b0000000_100101111110;
      15'b010_110101110110 : VALUE=19'b0000000_100101111110;
      15'b010_110101110111 : VALUE=19'b0000000_100101111110;
      15'b010_110101111000 : VALUE=19'b0000000_100101111110;
      15'b010_110101111001 : VALUE=19'b0000000_100101111110;
      15'b010_110101111010 : VALUE=19'b0000000_100101111110;
      15'b010_110101111011 : VALUE=19'b0000000_100101111101;
      15'b010_110101111100 : VALUE=19'b0000000_100101111101;
      15'b010_110101111101 : VALUE=19'b0000000_100101111101;
      15'b010_110101111110 : VALUE=19'b0000000_100101111101;
      15'b010_110101111111 : VALUE=19'b0000000_100101111101;
      15'b010_110110000000 : VALUE=19'b0000000_100101111101;
      15'b010_110110000001 : VALUE=19'b0000000_100101111101;
      15'b010_110110000010 : VALUE=19'b0000000_100101111101;
      15'b010_110110000011 : VALUE=19'b0000000_100101111101;
      15'b010_110110000100 : VALUE=19'b0000000_100101111101;
      15'b010_110110000101 : VALUE=19'b0000000_100101111100;
      15'b010_110110000110 : VALUE=19'b0000000_100101111100;
      15'b010_110110000111 : VALUE=19'b0000000_100101111100;
      15'b010_110110001000 : VALUE=19'b0000000_100101111100;
      15'b010_110110001001 : VALUE=19'b0000000_100101111100;
      15'b010_110110001010 : VALUE=19'b0000000_100101111100;
      15'b010_110110001011 : VALUE=19'b0000000_100101111100;
      15'b010_110110001100 : VALUE=19'b0000000_100101111100;
      15'b010_110110001101 : VALUE=19'b0000000_100101111100;
      15'b010_110110001110 : VALUE=19'b0000000_100101111011;
      15'b010_110110001111 : VALUE=19'b0000000_100101111011;
      15'b010_110110010000 : VALUE=19'b0000000_100101111011;
      15'b010_110110010001 : VALUE=19'b0000000_100101111011;
      15'b010_110110010010 : VALUE=19'b0000000_100101111011;
      15'b010_110110010011 : VALUE=19'b0000000_100101111011;
      15'b010_110110010100 : VALUE=19'b0000000_100101111011;
      15'b010_110110010101 : VALUE=19'b0000000_100101111011;
      15'b010_110110010110 : VALUE=19'b0000000_100101111011;
      15'b010_110110010111 : VALUE=19'b0000000_100101111011;
      15'b010_110110011000 : VALUE=19'b0000000_100101111010;
      15'b010_110110011001 : VALUE=19'b0000000_100101111010;
      15'b010_110110011010 : VALUE=19'b0000000_100101111010;
      15'b010_110110011011 : VALUE=19'b0000000_100101111010;
      15'b010_110110011100 : VALUE=19'b0000000_100101111010;
      15'b010_110110011101 : VALUE=19'b0000000_100101111010;
      15'b010_110110011110 : VALUE=19'b0000000_100101111010;
      15'b010_110110011111 : VALUE=19'b0000000_100101111010;
      15'b010_110110100000 : VALUE=19'b0000000_100101111010;
      15'b010_110110100001 : VALUE=19'b0000000_100101111001;
      15'b010_110110100010 : VALUE=19'b0000000_100101111001;
      15'b010_110110100011 : VALUE=19'b0000000_100101111001;
      15'b010_110110100100 : VALUE=19'b0000000_100101111001;
      15'b010_110110100101 : VALUE=19'b0000000_100101111001;
      15'b010_110110100110 : VALUE=19'b0000000_100101111001;
      15'b010_110110100111 : VALUE=19'b0000000_100101111001;
      15'b010_110110101000 : VALUE=19'b0000000_100101111001;
      15'b010_110110101001 : VALUE=19'b0000000_100101111001;
      15'b010_110110101010 : VALUE=19'b0000000_100101111001;
      15'b010_110110101011 : VALUE=19'b0000000_100101111000;
      15'b010_110110101100 : VALUE=19'b0000000_100101111000;
      15'b010_110110101101 : VALUE=19'b0000000_100101111000;
      15'b010_110110101110 : VALUE=19'b0000000_100101111000;
      15'b010_110110101111 : VALUE=19'b0000000_100101111000;
      15'b010_110110110000 : VALUE=19'b0000000_100101111000;
      15'b010_110110110001 : VALUE=19'b0000000_100101111000;
      15'b010_110110110010 : VALUE=19'b0000000_100101111000;
      15'b010_110110110011 : VALUE=19'b0000000_100101111000;
      15'b010_110110110100 : VALUE=19'b0000000_100101111000;
      15'b010_110110110101 : VALUE=19'b0000000_100101110111;
      15'b010_110110110110 : VALUE=19'b0000000_100101110111;
      15'b010_110110110111 : VALUE=19'b0000000_100101110111;
      15'b010_110110111000 : VALUE=19'b0000000_100101110111;
      15'b010_110110111001 : VALUE=19'b0000000_100101110111;
      15'b010_110110111010 : VALUE=19'b0000000_100101110111;
      15'b010_110110111011 : VALUE=19'b0000000_100101110111;
      15'b010_110110111100 : VALUE=19'b0000000_100101110111;
      15'b010_110110111101 : VALUE=19'b0000000_100101110111;
      15'b010_110110111110 : VALUE=19'b0000000_100101110110;
      15'b010_110110111111 : VALUE=19'b0000000_100101110110;
      15'b010_110111000000 : VALUE=19'b0000000_100101110110;
      15'b010_110111000001 : VALUE=19'b0000000_100101110110;
      15'b010_110111000010 : VALUE=19'b0000000_100101110110;
      15'b010_110111000011 : VALUE=19'b0000000_100101110110;
      15'b010_110111000100 : VALUE=19'b0000000_100101110110;
      15'b010_110111000101 : VALUE=19'b0000000_100101110110;
      15'b010_110111000110 : VALUE=19'b0000000_100101110110;
      15'b010_110111000111 : VALUE=19'b0000000_100101110110;
      15'b010_110111001000 : VALUE=19'b0000000_100101110101;
      15'b010_110111001001 : VALUE=19'b0000000_100101110101;
      15'b010_110111001010 : VALUE=19'b0000000_100101110101;
      15'b010_110111001011 : VALUE=19'b0000000_100101110101;
      15'b010_110111001100 : VALUE=19'b0000000_100101110101;
      15'b010_110111001101 : VALUE=19'b0000000_100101110101;
      15'b010_110111001110 : VALUE=19'b0000000_100101110101;
      15'b010_110111001111 : VALUE=19'b0000000_100101110101;
      15'b010_110111010000 : VALUE=19'b0000000_100101110101;
      15'b010_110111010001 : VALUE=19'b0000000_100101110101;
      15'b010_110111010010 : VALUE=19'b0000000_100101110100;
      15'b010_110111010011 : VALUE=19'b0000000_100101110100;
      15'b010_110111010100 : VALUE=19'b0000000_100101110100;
      15'b010_110111010101 : VALUE=19'b0000000_100101110100;
      15'b010_110111010110 : VALUE=19'b0000000_100101110100;
      15'b010_110111010111 : VALUE=19'b0000000_100101110100;
      15'b010_110111011000 : VALUE=19'b0000000_100101110100;
      15'b010_110111011001 : VALUE=19'b0000000_100101110100;
      15'b010_110111011010 : VALUE=19'b0000000_100101110100;
      15'b010_110111011011 : VALUE=19'b0000000_100101110011;
      15'b010_110111011100 : VALUE=19'b0000000_100101110011;
      15'b010_110111011101 : VALUE=19'b0000000_100101110011;
      15'b010_110111011110 : VALUE=19'b0000000_100101110011;
      15'b010_110111011111 : VALUE=19'b0000000_100101110011;
      15'b010_110111100000 : VALUE=19'b0000000_100101110011;
      15'b010_110111100001 : VALUE=19'b0000000_100101110011;
      15'b010_110111100010 : VALUE=19'b0000000_100101110011;
      15'b010_110111100011 : VALUE=19'b0000000_100101110011;
      15'b010_110111100100 : VALUE=19'b0000000_100101110011;
      15'b010_110111100101 : VALUE=19'b0000000_100101110010;
      15'b010_110111100110 : VALUE=19'b0000000_100101110010;
      15'b010_110111100111 : VALUE=19'b0000000_100101110010;
      15'b010_110111101000 : VALUE=19'b0000000_100101110010;
      15'b010_110111101001 : VALUE=19'b0000000_100101110010;
      15'b010_110111101010 : VALUE=19'b0000000_100101110010;
      15'b010_110111101011 : VALUE=19'b0000000_100101110010;
      15'b010_110111101100 : VALUE=19'b0000000_100101110010;
      15'b010_110111101101 : VALUE=19'b0000000_100101110010;
      15'b010_110111101110 : VALUE=19'b0000000_100101110010;
      15'b010_110111101111 : VALUE=19'b0000000_100101110001;
      15'b010_110111110000 : VALUE=19'b0000000_100101110001;
      15'b010_110111110001 : VALUE=19'b0000000_100101110001;
      15'b010_110111110010 : VALUE=19'b0000000_100101110001;
      15'b010_110111110011 : VALUE=19'b0000000_100101110001;
      15'b010_110111110100 : VALUE=19'b0000000_100101110001;
      15'b010_110111110101 : VALUE=19'b0000000_100101110001;
      15'b010_110111110110 : VALUE=19'b0000000_100101110001;
      15'b010_110111110111 : VALUE=19'b0000000_100101110001;
      15'b010_110111111000 : VALUE=19'b0000000_100101110001;
      15'b010_110111111001 : VALUE=19'b0000000_100101110000;
      15'b010_110111111010 : VALUE=19'b0000000_100101110000;
      15'b010_110111111011 : VALUE=19'b0000000_100101110000;
      15'b010_110111111100 : VALUE=19'b0000000_100101110000;
      15'b010_110111111101 : VALUE=19'b0000000_100101110000;
      15'b010_110111111110 : VALUE=19'b0000000_100101110000;
      15'b010_110111111111 : VALUE=19'b0000000_100101110000;
      15'b010_111000000000 : VALUE=19'b0000000_100101110000;
      15'b010_111000000001 : VALUE=19'b0000000_100101110000;
      15'b010_111000000010 : VALUE=19'b0000000_100101101111;
      15'b010_111000000011 : VALUE=19'b0000000_100101101111;
      15'b010_111000000100 : VALUE=19'b0000000_100101101111;
      15'b010_111000000101 : VALUE=19'b0000000_100101101111;
      15'b010_111000000110 : VALUE=19'b0000000_100101101111;
      15'b010_111000000111 : VALUE=19'b0000000_100101101111;
      15'b010_111000001000 : VALUE=19'b0000000_100101101111;
      15'b010_111000001001 : VALUE=19'b0000000_100101101111;
      15'b010_111000001010 : VALUE=19'b0000000_100101101111;
      15'b010_111000001011 : VALUE=19'b0000000_100101101111;
      15'b010_111000001100 : VALUE=19'b0000000_100101101110;
      15'b010_111000001101 : VALUE=19'b0000000_100101101110;
      15'b010_111000001110 : VALUE=19'b0000000_100101101110;
      15'b010_111000001111 : VALUE=19'b0000000_100101101110;
      15'b010_111000010000 : VALUE=19'b0000000_100101101110;
      15'b010_111000010001 : VALUE=19'b0000000_100101101110;
      15'b010_111000010010 : VALUE=19'b0000000_100101101110;
      15'b010_111000010011 : VALUE=19'b0000000_100101101110;
      15'b010_111000010100 : VALUE=19'b0000000_100101101110;
      15'b010_111000010101 : VALUE=19'b0000000_100101101110;
      15'b010_111000010110 : VALUE=19'b0000000_100101101101;
      15'b010_111000010111 : VALUE=19'b0000000_100101101101;
      15'b010_111000011000 : VALUE=19'b0000000_100101101101;
      15'b010_111000011001 : VALUE=19'b0000000_100101101101;
      15'b010_111000011010 : VALUE=19'b0000000_100101101101;
      15'b010_111000011011 : VALUE=19'b0000000_100101101101;
      15'b010_111000011100 : VALUE=19'b0000000_100101101101;
      15'b010_111000011101 : VALUE=19'b0000000_100101101101;
      15'b010_111000011110 : VALUE=19'b0000000_100101101101;
      15'b010_111000011111 : VALUE=19'b0000000_100101101101;
      15'b010_111000100000 : VALUE=19'b0000000_100101101100;
      15'b010_111000100001 : VALUE=19'b0000000_100101101100;
      15'b010_111000100010 : VALUE=19'b0000000_100101101100;
      15'b010_111000100011 : VALUE=19'b0000000_100101101100;
      15'b010_111000100100 : VALUE=19'b0000000_100101101100;
      15'b010_111000100101 : VALUE=19'b0000000_100101101100;
      15'b010_111000100110 : VALUE=19'b0000000_100101101100;
      15'b010_111000100111 : VALUE=19'b0000000_100101101100;
      15'b010_111000101000 : VALUE=19'b0000000_100101101100;
      15'b010_111000101001 : VALUE=19'b0000000_100101101011;
      15'b010_111000101010 : VALUE=19'b0000000_100101101011;
      15'b010_111000101011 : VALUE=19'b0000000_100101101011;
      15'b010_111000101100 : VALUE=19'b0000000_100101101011;
      15'b010_111000101101 : VALUE=19'b0000000_100101101011;
      15'b010_111000101110 : VALUE=19'b0000000_100101101011;
      15'b010_111000101111 : VALUE=19'b0000000_100101101011;
      15'b010_111000110000 : VALUE=19'b0000000_100101101011;
      15'b010_111000110001 : VALUE=19'b0000000_100101101011;
      15'b010_111000110010 : VALUE=19'b0000000_100101101011;
      15'b010_111000110011 : VALUE=19'b0000000_100101101010;
      15'b010_111000110100 : VALUE=19'b0000000_100101101010;
      15'b010_111000110101 : VALUE=19'b0000000_100101101010;
      15'b010_111000110110 : VALUE=19'b0000000_100101101010;
      15'b010_111000110111 : VALUE=19'b0000000_100101101010;
      15'b010_111000111000 : VALUE=19'b0000000_100101101010;
      15'b010_111000111001 : VALUE=19'b0000000_100101101010;
      15'b010_111000111010 : VALUE=19'b0000000_100101101010;
      15'b010_111000111011 : VALUE=19'b0000000_100101101010;
      15'b010_111000111100 : VALUE=19'b0000000_100101101010;
      15'b010_111000111101 : VALUE=19'b0000000_100101101001;
      15'b010_111000111110 : VALUE=19'b0000000_100101101001;
      15'b010_111000111111 : VALUE=19'b0000000_100101101001;
      15'b010_111001000000 : VALUE=19'b0000000_100101101001;
      15'b010_111001000001 : VALUE=19'b0000000_100101101001;
      15'b010_111001000010 : VALUE=19'b0000000_100101101001;
      15'b010_111001000011 : VALUE=19'b0000000_100101101001;
      15'b010_111001000100 : VALUE=19'b0000000_100101101001;
      15'b010_111001000101 : VALUE=19'b0000000_100101101001;
      15'b010_111001000110 : VALUE=19'b0000000_100101101001;
      15'b010_111001000111 : VALUE=19'b0000000_100101101000;
      15'b010_111001001000 : VALUE=19'b0000000_100101101000;
      15'b010_111001001001 : VALUE=19'b0000000_100101101000;
      15'b010_111001001010 : VALUE=19'b0000000_100101101000;
      15'b010_111001001011 : VALUE=19'b0000000_100101101000;
      15'b010_111001001100 : VALUE=19'b0000000_100101101000;
      15'b010_111001001101 : VALUE=19'b0000000_100101101000;
      15'b010_111001001110 : VALUE=19'b0000000_100101101000;
      15'b010_111001001111 : VALUE=19'b0000000_100101101000;
      15'b010_111001010000 : VALUE=19'b0000000_100101101000;
      15'b010_111001010001 : VALUE=19'b0000000_100101100111;
      15'b010_111001010010 : VALUE=19'b0000000_100101100111;
      15'b010_111001010011 : VALUE=19'b0000000_100101100111;
      15'b010_111001010100 : VALUE=19'b0000000_100101100111;
      15'b010_111001010101 : VALUE=19'b0000000_100101100111;
      15'b010_111001010110 : VALUE=19'b0000000_100101100111;
      15'b010_111001010111 : VALUE=19'b0000000_100101100111;
      15'b010_111001011000 : VALUE=19'b0000000_100101100111;
      15'b010_111001011001 : VALUE=19'b0000000_100101100111;
      15'b010_111001011010 : VALUE=19'b0000000_100101100111;
      15'b010_111001011011 : VALUE=19'b0000000_100101100110;
      15'b010_111001011100 : VALUE=19'b0000000_100101100110;
      15'b010_111001011101 : VALUE=19'b0000000_100101100110;
      15'b010_111001011110 : VALUE=19'b0000000_100101100110;
      15'b010_111001011111 : VALUE=19'b0000000_100101100110;
      15'b010_111001100000 : VALUE=19'b0000000_100101100110;
      15'b010_111001100001 : VALUE=19'b0000000_100101100110;
      15'b010_111001100010 : VALUE=19'b0000000_100101100110;
      15'b010_111001100011 : VALUE=19'b0000000_100101100110;
      15'b010_111001100100 : VALUE=19'b0000000_100101100101;
      15'b010_111001100101 : VALUE=19'b0000000_100101100101;
      15'b010_111001100110 : VALUE=19'b0000000_100101100101;
      15'b010_111001100111 : VALUE=19'b0000000_100101100101;
      15'b010_111001101000 : VALUE=19'b0000000_100101100101;
      15'b010_111001101001 : VALUE=19'b0000000_100101100101;
      15'b010_111001101010 : VALUE=19'b0000000_100101100101;
      15'b010_111001101011 : VALUE=19'b0000000_100101100101;
      15'b010_111001101100 : VALUE=19'b0000000_100101100101;
      15'b010_111001101101 : VALUE=19'b0000000_100101100101;
      15'b010_111001101110 : VALUE=19'b0000000_100101100100;
      15'b010_111001101111 : VALUE=19'b0000000_100101100100;
      15'b010_111001110000 : VALUE=19'b0000000_100101100100;
      15'b010_111001110001 : VALUE=19'b0000000_100101100100;
      15'b010_111001110010 : VALUE=19'b0000000_100101100100;
      15'b010_111001110011 : VALUE=19'b0000000_100101100100;
      15'b010_111001110100 : VALUE=19'b0000000_100101100100;
      15'b010_111001110101 : VALUE=19'b0000000_100101100100;
      15'b010_111001110110 : VALUE=19'b0000000_100101100100;
      15'b010_111001110111 : VALUE=19'b0000000_100101100100;
      15'b010_111001111000 : VALUE=19'b0000000_100101100011;
      15'b010_111001111001 : VALUE=19'b0000000_100101100011;
      15'b010_111001111010 : VALUE=19'b0000000_100101100011;
      15'b010_111001111011 : VALUE=19'b0000000_100101100011;
      15'b010_111001111100 : VALUE=19'b0000000_100101100011;
      15'b010_111001111101 : VALUE=19'b0000000_100101100011;
      15'b010_111001111110 : VALUE=19'b0000000_100101100011;
      15'b010_111001111111 : VALUE=19'b0000000_100101100011;
      15'b010_111010000000 : VALUE=19'b0000000_100101100011;
      15'b010_111010000001 : VALUE=19'b0000000_100101100011;
      15'b010_111010000010 : VALUE=19'b0000000_100101100010;
      15'b010_111010000011 : VALUE=19'b0000000_100101100010;
      15'b010_111010000100 : VALUE=19'b0000000_100101100010;
      15'b010_111010000101 : VALUE=19'b0000000_100101100010;
      15'b010_111010000110 : VALUE=19'b0000000_100101100010;
      15'b010_111010000111 : VALUE=19'b0000000_100101100010;
      15'b010_111010001000 : VALUE=19'b0000000_100101100010;
      15'b010_111010001001 : VALUE=19'b0000000_100101100010;
      15'b010_111010001010 : VALUE=19'b0000000_100101100010;
      15'b010_111010001011 : VALUE=19'b0000000_100101100010;
      15'b010_111010001100 : VALUE=19'b0000000_100101100001;
      15'b010_111010001101 : VALUE=19'b0000000_100101100001;
      15'b010_111010001110 : VALUE=19'b0000000_100101100001;
      15'b010_111010001111 : VALUE=19'b0000000_100101100001;
      15'b010_111010010000 : VALUE=19'b0000000_100101100001;
      15'b010_111010010001 : VALUE=19'b0000000_100101100001;
      15'b010_111010010010 : VALUE=19'b0000000_100101100001;
      15'b010_111010010011 : VALUE=19'b0000000_100101100001;
      15'b010_111010010100 : VALUE=19'b0000000_100101100001;
      15'b010_111010010101 : VALUE=19'b0000000_100101100001;
      15'b010_111010010110 : VALUE=19'b0000000_100101100000;
      15'b010_111010010111 : VALUE=19'b0000000_100101100000;
      15'b010_111010011000 : VALUE=19'b0000000_100101100000;
      15'b010_111010011001 : VALUE=19'b0000000_100101100000;
      15'b010_111010011010 : VALUE=19'b0000000_100101100000;
      15'b010_111010011011 : VALUE=19'b0000000_100101100000;
      15'b010_111010011100 : VALUE=19'b0000000_100101100000;
      15'b010_111010011101 : VALUE=19'b0000000_100101100000;
      15'b010_111010011110 : VALUE=19'b0000000_100101100000;
      15'b010_111010011111 : VALUE=19'b0000000_100101100000;
      15'b010_111010100000 : VALUE=19'b0000000_100101011111;
      15'b010_111010100001 : VALUE=19'b0000000_100101011111;
      15'b010_111010100010 : VALUE=19'b0000000_100101011111;
      15'b010_111010100011 : VALUE=19'b0000000_100101011111;
      15'b010_111010100100 : VALUE=19'b0000000_100101011111;
      15'b010_111010100101 : VALUE=19'b0000000_100101011111;
      15'b010_111010100110 : VALUE=19'b0000000_100101011111;
      15'b010_111010100111 : VALUE=19'b0000000_100101011111;
      15'b010_111010101000 : VALUE=19'b0000000_100101011111;
      15'b010_111010101001 : VALUE=19'b0000000_100101011111;
      15'b010_111010101010 : VALUE=19'b0000000_100101011110;
      15'b010_111010101011 : VALUE=19'b0000000_100101011110;
      15'b010_111010101100 : VALUE=19'b0000000_100101011110;
      15'b010_111010101101 : VALUE=19'b0000000_100101011110;
      15'b010_111010101110 : VALUE=19'b0000000_100101011110;
      15'b010_111010101111 : VALUE=19'b0000000_100101011110;
      15'b010_111010110000 : VALUE=19'b0000000_100101011110;
      15'b010_111010110001 : VALUE=19'b0000000_100101011110;
      15'b010_111010110010 : VALUE=19'b0000000_100101011110;
      15'b010_111010110011 : VALUE=19'b0000000_100101011110;
      15'b010_111010110100 : VALUE=19'b0000000_100101011101;
      15'b010_111010110101 : VALUE=19'b0000000_100101011101;
      15'b010_111010110110 : VALUE=19'b0000000_100101011101;
      15'b010_111010110111 : VALUE=19'b0000000_100101011101;
      15'b010_111010111000 : VALUE=19'b0000000_100101011101;
      15'b010_111010111001 : VALUE=19'b0000000_100101011101;
      15'b010_111010111010 : VALUE=19'b0000000_100101011101;
      15'b010_111010111011 : VALUE=19'b0000000_100101011101;
      15'b010_111010111100 : VALUE=19'b0000000_100101011101;
      15'b010_111010111101 : VALUE=19'b0000000_100101011101;
      15'b010_111010111110 : VALUE=19'b0000000_100101011100;
      15'b010_111010111111 : VALUE=19'b0000000_100101011100;
      15'b010_111011000000 : VALUE=19'b0000000_100101011100;
      15'b010_111011000001 : VALUE=19'b0000000_100101011100;
      15'b010_111011000010 : VALUE=19'b0000000_100101011100;
      15'b010_111011000011 : VALUE=19'b0000000_100101011100;
      15'b010_111011000100 : VALUE=19'b0000000_100101011100;
      15'b010_111011000101 : VALUE=19'b0000000_100101011100;
      15'b010_111011000110 : VALUE=19'b0000000_100101011100;
      15'b010_111011000111 : VALUE=19'b0000000_100101011100;
      15'b010_111011001000 : VALUE=19'b0000000_100101011011;
      15'b010_111011001001 : VALUE=19'b0000000_100101011011;
      15'b010_111011001010 : VALUE=19'b0000000_100101011011;
      15'b010_111011001011 : VALUE=19'b0000000_100101011011;
      15'b010_111011001100 : VALUE=19'b0000000_100101011011;
      15'b010_111011001101 : VALUE=19'b0000000_100101011011;
      15'b010_111011001110 : VALUE=19'b0000000_100101011011;
      15'b010_111011001111 : VALUE=19'b0000000_100101011011;
      15'b010_111011010000 : VALUE=19'b0000000_100101011011;
      15'b010_111011010001 : VALUE=19'b0000000_100101011011;
      15'b010_111011010010 : VALUE=19'b0000000_100101011010;
      15'b010_111011010011 : VALUE=19'b0000000_100101011010;
      15'b010_111011010100 : VALUE=19'b0000000_100101011010;
      15'b010_111011010101 : VALUE=19'b0000000_100101011010;
      15'b010_111011010110 : VALUE=19'b0000000_100101011010;
      15'b010_111011010111 : VALUE=19'b0000000_100101011010;
      15'b010_111011011000 : VALUE=19'b0000000_100101011010;
      15'b010_111011011001 : VALUE=19'b0000000_100101011010;
      15'b010_111011011010 : VALUE=19'b0000000_100101011010;
      15'b010_111011011011 : VALUE=19'b0000000_100101011010;
      15'b010_111011011100 : VALUE=19'b0000000_100101011001;
      15'b010_111011011101 : VALUE=19'b0000000_100101011001;
      15'b010_111011011110 : VALUE=19'b0000000_100101011001;
      15'b010_111011011111 : VALUE=19'b0000000_100101011001;
      15'b010_111011100000 : VALUE=19'b0000000_100101011001;
      15'b010_111011100001 : VALUE=19'b0000000_100101011001;
      15'b010_111011100010 : VALUE=19'b0000000_100101011001;
      15'b010_111011100011 : VALUE=19'b0000000_100101011001;
      15'b010_111011100100 : VALUE=19'b0000000_100101011001;
      15'b010_111011100101 : VALUE=19'b0000000_100101011001;
      15'b010_111011100110 : VALUE=19'b0000000_100101011000;
      15'b010_111011100111 : VALUE=19'b0000000_100101011000;
      15'b010_111011101000 : VALUE=19'b0000000_100101011000;
      15'b010_111011101001 : VALUE=19'b0000000_100101011000;
      15'b010_111011101010 : VALUE=19'b0000000_100101011000;
      15'b010_111011101011 : VALUE=19'b0000000_100101011000;
      15'b010_111011101100 : VALUE=19'b0000000_100101011000;
      15'b010_111011101101 : VALUE=19'b0000000_100101011000;
      15'b010_111011101110 : VALUE=19'b0000000_100101011000;
      15'b010_111011101111 : VALUE=19'b0000000_100101011000;
      15'b010_111011110000 : VALUE=19'b0000000_100101010111;
      15'b010_111011110001 : VALUE=19'b0000000_100101010111;
      15'b010_111011110010 : VALUE=19'b0000000_100101010111;
      15'b010_111011110011 : VALUE=19'b0000000_100101010111;
      15'b010_111011110100 : VALUE=19'b0000000_100101010111;
      15'b010_111011110101 : VALUE=19'b0000000_100101010111;
      15'b010_111011110110 : VALUE=19'b0000000_100101010111;
      15'b010_111011110111 : VALUE=19'b0000000_100101010111;
      15'b010_111011111000 : VALUE=19'b0000000_100101010111;
      15'b010_111011111001 : VALUE=19'b0000000_100101010111;
      15'b010_111011111010 : VALUE=19'b0000000_100101010110;
      15'b010_111011111011 : VALUE=19'b0000000_100101010110;
      15'b010_111011111100 : VALUE=19'b0000000_100101010110;
      15'b010_111011111101 : VALUE=19'b0000000_100101010110;
      15'b010_111011111110 : VALUE=19'b0000000_100101010110;
      15'b010_111011111111 : VALUE=19'b0000000_100101010110;
      15'b010_111100000000 : VALUE=19'b0000000_100101010110;
      15'b010_111100000001 : VALUE=19'b0000000_100101010110;
      15'b010_111100000010 : VALUE=19'b0000000_100101010110;
      15'b010_111100000011 : VALUE=19'b0000000_100101010110;
      15'b010_111100000100 : VALUE=19'b0000000_100101010101;
      15'b010_111100000101 : VALUE=19'b0000000_100101010101;
      15'b010_111100000110 : VALUE=19'b0000000_100101010101;
      15'b010_111100000111 : VALUE=19'b0000000_100101010101;
      15'b010_111100001000 : VALUE=19'b0000000_100101010101;
      15'b010_111100001001 : VALUE=19'b0000000_100101010101;
      15'b010_111100001010 : VALUE=19'b0000000_100101010101;
      15'b010_111100001011 : VALUE=19'b0000000_100101010101;
      15'b010_111100001100 : VALUE=19'b0000000_100101010101;
      15'b010_111100001101 : VALUE=19'b0000000_100101010101;
      15'b010_111100001110 : VALUE=19'b0000000_100101010100;
      15'b010_111100001111 : VALUE=19'b0000000_100101010100;
      15'b010_111100010000 : VALUE=19'b0000000_100101010100;
      15'b010_111100010001 : VALUE=19'b0000000_100101010100;
      15'b010_111100010010 : VALUE=19'b0000000_100101010100;
      15'b010_111100010011 : VALUE=19'b0000000_100101010100;
      15'b010_111100010100 : VALUE=19'b0000000_100101010100;
      15'b010_111100010101 : VALUE=19'b0000000_100101010100;
      15'b010_111100010110 : VALUE=19'b0000000_100101010100;
      15'b010_111100010111 : VALUE=19'b0000000_100101010100;
      15'b010_111100011000 : VALUE=19'b0000000_100101010011;
      15'b010_111100011001 : VALUE=19'b0000000_100101010011;
      15'b010_111100011010 : VALUE=19'b0000000_100101010011;
      15'b010_111100011011 : VALUE=19'b0000000_100101010011;
      15'b010_111100011100 : VALUE=19'b0000000_100101010011;
      15'b010_111100011101 : VALUE=19'b0000000_100101010011;
      15'b010_111100011110 : VALUE=19'b0000000_100101010011;
      15'b010_111100011111 : VALUE=19'b0000000_100101010011;
      15'b010_111100100000 : VALUE=19'b0000000_100101010011;
      15'b010_111100100001 : VALUE=19'b0000000_100101010011;
      15'b010_111100100010 : VALUE=19'b0000000_100101010010;
      15'b010_111100100011 : VALUE=19'b0000000_100101010010;
      15'b010_111100100100 : VALUE=19'b0000000_100101010010;
      15'b010_111100100101 : VALUE=19'b0000000_100101010010;
      15'b010_111100100110 : VALUE=19'b0000000_100101010010;
      15'b010_111100100111 : VALUE=19'b0000000_100101010010;
      15'b010_111100101000 : VALUE=19'b0000000_100101010010;
      15'b010_111100101001 : VALUE=19'b0000000_100101010010;
      15'b010_111100101010 : VALUE=19'b0000000_100101010010;
      15'b010_111100101011 : VALUE=19'b0000000_100101010010;
      15'b010_111100101100 : VALUE=19'b0000000_100101010001;
      15'b010_111100101101 : VALUE=19'b0000000_100101010001;
      15'b010_111100101110 : VALUE=19'b0000000_100101010001;
      15'b010_111100101111 : VALUE=19'b0000000_100101010001;
      15'b010_111100110000 : VALUE=19'b0000000_100101010001;
      15'b010_111100110001 : VALUE=19'b0000000_100101010001;
      15'b010_111100110010 : VALUE=19'b0000000_100101010001;
      15'b010_111100110011 : VALUE=19'b0000000_100101010001;
      15'b010_111100110100 : VALUE=19'b0000000_100101010001;
      15'b010_111100110101 : VALUE=19'b0000000_100101010001;
      15'b010_111100110110 : VALUE=19'b0000000_100101010001;
      15'b010_111100110111 : VALUE=19'b0000000_100101010000;
      15'b010_111100111000 : VALUE=19'b0000000_100101010000;
      15'b010_111100111001 : VALUE=19'b0000000_100101010000;
      15'b010_111100111010 : VALUE=19'b0000000_100101010000;
      15'b010_111100111011 : VALUE=19'b0000000_100101010000;
      15'b010_111100111100 : VALUE=19'b0000000_100101010000;
      15'b010_111100111101 : VALUE=19'b0000000_100101010000;
      15'b010_111100111110 : VALUE=19'b0000000_100101010000;
      15'b010_111100111111 : VALUE=19'b0000000_100101010000;
      15'b010_111101000000 : VALUE=19'b0000000_100101010000;
      15'b010_111101000001 : VALUE=19'b0000000_100101001111;
      15'b010_111101000010 : VALUE=19'b0000000_100101001111;
      15'b010_111101000011 : VALUE=19'b0000000_100101001111;
      15'b010_111101000100 : VALUE=19'b0000000_100101001111;
      15'b010_111101000101 : VALUE=19'b0000000_100101001111;
      15'b010_111101000110 : VALUE=19'b0000000_100101001111;
      15'b010_111101000111 : VALUE=19'b0000000_100101001111;
      15'b010_111101001000 : VALUE=19'b0000000_100101001111;
      15'b010_111101001001 : VALUE=19'b0000000_100101001111;
      15'b010_111101001010 : VALUE=19'b0000000_100101001111;
      15'b010_111101001011 : VALUE=19'b0000000_100101001110;
      15'b010_111101001100 : VALUE=19'b0000000_100101001110;
      15'b010_111101001101 : VALUE=19'b0000000_100101001110;
      15'b010_111101001110 : VALUE=19'b0000000_100101001110;
      15'b010_111101001111 : VALUE=19'b0000000_100101001110;
      15'b010_111101010000 : VALUE=19'b0000000_100101001110;
      15'b010_111101010001 : VALUE=19'b0000000_100101001110;
      15'b010_111101010010 : VALUE=19'b0000000_100101001110;
      15'b010_111101010011 : VALUE=19'b0000000_100101001110;
      15'b010_111101010100 : VALUE=19'b0000000_100101001110;
      15'b010_111101010101 : VALUE=19'b0000000_100101001101;
      15'b010_111101010110 : VALUE=19'b0000000_100101001101;
      15'b010_111101010111 : VALUE=19'b0000000_100101001101;
      15'b010_111101011000 : VALUE=19'b0000000_100101001101;
      15'b010_111101011001 : VALUE=19'b0000000_100101001101;
      15'b010_111101011010 : VALUE=19'b0000000_100101001101;
      15'b010_111101011011 : VALUE=19'b0000000_100101001101;
      15'b010_111101011100 : VALUE=19'b0000000_100101001101;
      15'b010_111101011101 : VALUE=19'b0000000_100101001101;
      15'b010_111101011110 : VALUE=19'b0000000_100101001101;
      15'b010_111101011111 : VALUE=19'b0000000_100101001100;
      15'b010_111101100000 : VALUE=19'b0000000_100101001100;
      15'b010_111101100001 : VALUE=19'b0000000_100101001100;
      15'b010_111101100010 : VALUE=19'b0000000_100101001100;
      15'b010_111101100011 : VALUE=19'b0000000_100101001100;
      15'b010_111101100100 : VALUE=19'b0000000_100101001100;
      15'b010_111101100101 : VALUE=19'b0000000_100101001100;
      15'b010_111101100110 : VALUE=19'b0000000_100101001100;
      15'b010_111101100111 : VALUE=19'b0000000_100101001100;
      15'b010_111101101000 : VALUE=19'b0000000_100101001100;
      15'b010_111101101001 : VALUE=19'b0000000_100101001011;
      15'b010_111101101010 : VALUE=19'b0000000_100101001011;
      15'b010_111101101011 : VALUE=19'b0000000_100101001011;
      15'b010_111101101100 : VALUE=19'b0000000_100101001011;
      15'b010_111101101101 : VALUE=19'b0000000_100101001011;
      15'b010_111101101110 : VALUE=19'b0000000_100101001011;
      15'b010_111101101111 : VALUE=19'b0000000_100101001011;
      15'b010_111101110000 : VALUE=19'b0000000_100101001011;
      15'b010_111101110001 : VALUE=19'b0000000_100101001011;
      15'b010_111101110010 : VALUE=19'b0000000_100101001011;
      15'b010_111101110011 : VALUE=19'b0000000_100101001011;
      15'b010_111101110100 : VALUE=19'b0000000_100101001010;
      15'b010_111101110101 : VALUE=19'b0000000_100101001010;
      15'b010_111101110110 : VALUE=19'b0000000_100101001010;
      15'b010_111101110111 : VALUE=19'b0000000_100101001010;
      15'b010_111101111000 : VALUE=19'b0000000_100101001010;
      15'b010_111101111001 : VALUE=19'b0000000_100101001010;
      15'b010_111101111010 : VALUE=19'b0000000_100101001010;
      15'b010_111101111011 : VALUE=19'b0000000_100101001010;
      15'b010_111101111100 : VALUE=19'b0000000_100101001010;
      15'b010_111101111101 : VALUE=19'b0000000_100101001010;
      15'b010_111101111110 : VALUE=19'b0000000_100101001001;
      15'b010_111101111111 : VALUE=19'b0000000_100101001001;
      15'b010_111110000000 : VALUE=19'b0000000_100101001001;
      15'b010_111110000001 : VALUE=19'b0000000_100101001001;
      15'b010_111110000010 : VALUE=19'b0000000_100101001001;
      15'b010_111110000011 : VALUE=19'b0000000_100101001001;
      15'b010_111110000100 : VALUE=19'b0000000_100101001001;
      15'b010_111110000101 : VALUE=19'b0000000_100101001001;
      15'b010_111110000110 : VALUE=19'b0000000_100101001001;
      15'b010_111110000111 : VALUE=19'b0000000_100101001001;
      15'b010_111110001000 : VALUE=19'b0000000_100101001000;
      15'b010_111110001001 : VALUE=19'b0000000_100101001000;
      15'b010_111110001010 : VALUE=19'b0000000_100101001000;
      15'b010_111110001011 : VALUE=19'b0000000_100101001000;
      15'b010_111110001100 : VALUE=19'b0000000_100101001000;
      15'b010_111110001101 : VALUE=19'b0000000_100101001000;
      15'b010_111110001110 : VALUE=19'b0000000_100101001000;
      15'b010_111110001111 : VALUE=19'b0000000_100101001000;
      15'b010_111110010000 : VALUE=19'b0000000_100101001000;
      15'b010_111110010001 : VALUE=19'b0000000_100101001000;
      15'b010_111110010010 : VALUE=19'b0000000_100101000111;
      15'b010_111110010011 : VALUE=19'b0000000_100101000111;
      15'b010_111110010100 : VALUE=19'b0000000_100101000111;
      15'b010_111110010101 : VALUE=19'b0000000_100101000111;
      15'b010_111110010110 : VALUE=19'b0000000_100101000111;
      15'b010_111110010111 : VALUE=19'b0000000_100101000111;
      15'b010_111110011000 : VALUE=19'b0000000_100101000111;
      15'b010_111110011001 : VALUE=19'b0000000_100101000111;
      15'b010_111110011010 : VALUE=19'b0000000_100101000111;
      15'b010_111110011011 : VALUE=19'b0000000_100101000111;
      15'b010_111110011100 : VALUE=19'b0000000_100101000111;
      15'b010_111110011101 : VALUE=19'b0000000_100101000110;
      15'b010_111110011110 : VALUE=19'b0000000_100101000110;
      15'b010_111110011111 : VALUE=19'b0000000_100101000110;
      15'b010_111110100000 : VALUE=19'b0000000_100101000110;
      15'b010_111110100001 : VALUE=19'b0000000_100101000110;
      15'b010_111110100010 : VALUE=19'b0000000_100101000110;
      15'b010_111110100011 : VALUE=19'b0000000_100101000110;
      15'b010_111110100100 : VALUE=19'b0000000_100101000110;
      15'b010_111110100101 : VALUE=19'b0000000_100101000110;
      15'b010_111110100110 : VALUE=19'b0000000_100101000110;
      15'b010_111110100111 : VALUE=19'b0000000_100101000101;
      15'b010_111110101000 : VALUE=19'b0000000_100101000101;
      15'b010_111110101001 : VALUE=19'b0000000_100101000101;
      15'b010_111110101010 : VALUE=19'b0000000_100101000101;
      15'b010_111110101011 : VALUE=19'b0000000_100101000101;
      15'b010_111110101100 : VALUE=19'b0000000_100101000101;
      15'b010_111110101101 : VALUE=19'b0000000_100101000101;
      15'b010_111110101110 : VALUE=19'b0000000_100101000101;
      15'b010_111110101111 : VALUE=19'b0000000_100101000101;
      15'b010_111110110000 : VALUE=19'b0000000_100101000101;
      15'b010_111110110001 : VALUE=19'b0000000_100101000100;
      15'b010_111110110010 : VALUE=19'b0000000_100101000100;
      15'b010_111110110011 : VALUE=19'b0000000_100101000100;
      15'b010_111110110100 : VALUE=19'b0000000_100101000100;
      15'b010_111110110101 : VALUE=19'b0000000_100101000100;
      15'b010_111110110110 : VALUE=19'b0000000_100101000100;
      15'b010_111110110111 : VALUE=19'b0000000_100101000100;
      15'b010_111110111000 : VALUE=19'b0000000_100101000100;
      15'b010_111110111001 : VALUE=19'b0000000_100101000100;
      15'b010_111110111010 : VALUE=19'b0000000_100101000100;
      15'b010_111110111011 : VALUE=19'b0000000_100101000011;
      15'b010_111110111100 : VALUE=19'b0000000_100101000011;
      15'b010_111110111101 : VALUE=19'b0000000_100101000011;
      15'b010_111110111110 : VALUE=19'b0000000_100101000011;
      15'b010_111110111111 : VALUE=19'b0000000_100101000011;
      15'b010_111111000000 : VALUE=19'b0000000_100101000011;
      15'b010_111111000001 : VALUE=19'b0000000_100101000011;
      15'b010_111111000010 : VALUE=19'b0000000_100101000011;
      15'b010_111111000011 : VALUE=19'b0000000_100101000011;
      15'b010_111111000100 : VALUE=19'b0000000_100101000011;
      15'b010_111111000101 : VALUE=19'b0000000_100101000011;
      15'b010_111111000110 : VALUE=19'b0000000_100101000010;
      15'b010_111111000111 : VALUE=19'b0000000_100101000010;
      15'b010_111111001000 : VALUE=19'b0000000_100101000010;
      15'b010_111111001001 : VALUE=19'b0000000_100101000010;
      15'b010_111111001010 : VALUE=19'b0000000_100101000010;
      15'b010_111111001011 : VALUE=19'b0000000_100101000010;
      15'b010_111111001100 : VALUE=19'b0000000_100101000010;
      15'b010_111111001101 : VALUE=19'b0000000_100101000010;
      15'b010_111111001110 : VALUE=19'b0000000_100101000010;
      15'b010_111111001111 : VALUE=19'b0000000_100101000010;
      15'b010_111111010000 : VALUE=19'b0000000_100101000001;
      15'b010_111111010001 : VALUE=19'b0000000_100101000001;
      15'b010_111111010010 : VALUE=19'b0000000_100101000001;
      15'b010_111111010011 : VALUE=19'b0000000_100101000001;
      15'b010_111111010100 : VALUE=19'b0000000_100101000001;
      15'b010_111111010101 : VALUE=19'b0000000_100101000001;
      15'b010_111111010110 : VALUE=19'b0000000_100101000001;
      15'b010_111111010111 : VALUE=19'b0000000_100101000001;
      15'b010_111111011000 : VALUE=19'b0000000_100101000001;
      15'b010_111111011001 : VALUE=19'b0000000_100101000001;
      15'b010_111111011010 : VALUE=19'b0000000_100101000000;
      15'b010_111111011011 : VALUE=19'b0000000_100101000000;
      15'b010_111111011100 : VALUE=19'b0000000_100101000000;
      15'b010_111111011101 : VALUE=19'b0000000_100101000000;
      15'b010_111111011110 : VALUE=19'b0000000_100101000000;
      15'b010_111111011111 : VALUE=19'b0000000_100101000000;
      15'b010_111111100000 : VALUE=19'b0000000_100101000000;
      15'b010_111111100001 : VALUE=19'b0000000_100101000000;
      15'b010_111111100010 : VALUE=19'b0000000_100101000000;
      15'b010_111111100011 : VALUE=19'b0000000_100101000000;
      15'b010_111111100100 : VALUE=19'b0000000_100101000000;
      15'b010_111111100101 : VALUE=19'b0000000_100100111111;
      15'b010_111111100110 : VALUE=19'b0000000_100100111111;
      15'b010_111111100111 : VALUE=19'b0000000_100100111111;
      15'b010_111111101000 : VALUE=19'b0000000_100100111111;
      15'b010_111111101001 : VALUE=19'b0000000_100100111111;
      15'b010_111111101010 : VALUE=19'b0000000_100100111111;
      15'b010_111111101011 : VALUE=19'b0000000_100100111111;
      15'b010_111111101100 : VALUE=19'b0000000_100100111111;
      15'b010_111111101101 : VALUE=19'b0000000_100100111111;
      15'b010_111111101110 : VALUE=19'b0000000_100100111111;
      15'b010_111111101111 : VALUE=19'b0000000_100100111110;
      15'b010_111111110000 : VALUE=19'b0000000_100100111110;
      15'b010_111111110001 : VALUE=19'b0000000_100100111110;
      15'b010_111111110010 : VALUE=19'b0000000_100100111110;
      15'b010_111111110011 : VALUE=19'b0000000_100100111110;
      15'b010_111111110100 : VALUE=19'b0000000_100100111110;
      15'b010_111111110101 : VALUE=19'b0000000_100100111110;
      15'b010_111111110110 : VALUE=19'b0000000_100100111110;
      15'b010_111111110111 : VALUE=19'b0000000_100100111110;
      15'b010_111111111000 : VALUE=19'b0000000_100100111110;
      15'b010_111111111001 : VALUE=19'b0000000_100100111110;
      15'b010_111111111010 : VALUE=19'b0000000_100100111101;
      15'b010_111111111011 : VALUE=19'b0000000_100100111101;
      15'b010_111111111100 : VALUE=19'b0000000_100100111101;
      15'b010_111111111101 : VALUE=19'b0000000_100100111101;
      15'b010_111111111110 : VALUE=19'b0000000_100100111101;
      15'b010_111111111111 : VALUE=19'b0000000_100100111101;
      15'b011_000000000000 : VALUE=19'b0000000_100100111101;
      15'b011_000000000001 : VALUE=19'b0000000_100100111101;
      15'b011_000000000010 : VALUE=19'b0000000_100100111101;
      15'b011_000000000011 : VALUE=19'b0000000_100100111101;
      15'b011_000000000100 : VALUE=19'b0000000_100100111100;
      15'b011_000000000101 : VALUE=19'b0000000_100100111100;
      15'b011_000000000110 : VALUE=19'b0000000_100100111100;
      15'b011_000000000111 : VALUE=19'b0000000_100100111100;
      15'b011_000000001000 : VALUE=19'b0000000_100100111100;
      15'b011_000000001001 : VALUE=19'b0000000_100100111100;
      15'b011_000000001010 : VALUE=19'b0000000_100100111100;
      15'b011_000000001011 : VALUE=19'b0000000_100100111100;
      15'b011_000000001100 : VALUE=19'b0000000_100100111100;
      15'b011_000000001101 : VALUE=19'b0000000_100100111100;
      15'b011_000000001110 : VALUE=19'b0000000_100100111011;
      15'b011_000000001111 : VALUE=19'b0000000_100100111011;
      15'b011_000000010000 : VALUE=19'b0000000_100100111011;
      15'b011_000000010001 : VALUE=19'b0000000_100100111011;
      15'b011_000000010010 : VALUE=19'b0000000_100100111011;
      15'b011_000000010011 : VALUE=19'b0000000_100100111011;
      15'b011_000000010100 : VALUE=19'b0000000_100100111011;
      15'b011_000000010101 : VALUE=19'b0000000_100100111011;
      15'b011_000000010110 : VALUE=19'b0000000_100100111011;
      15'b011_000000010111 : VALUE=19'b0000000_100100111011;
      15'b011_000000011000 : VALUE=19'b0000000_100100111011;
      15'b011_000000011001 : VALUE=19'b0000000_100100111010;
      15'b011_000000011010 : VALUE=19'b0000000_100100111010;
      15'b011_000000011011 : VALUE=19'b0000000_100100111010;
      15'b011_000000011100 : VALUE=19'b0000000_100100111010;
      15'b011_000000011101 : VALUE=19'b0000000_100100111010;
      15'b011_000000011110 : VALUE=19'b0000000_100100111010;
      15'b011_000000011111 : VALUE=19'b0000000_100100111010;
      15'b011_000000100000 : VALUE=19'b0000000_100100111010;
      15'b011_000000100001 : VALUE=19'b0000000_100100111010;
      15'b011_000000100010 : VALUE=19'b0000000_100100111010;
      15'b011_000000100011 : VALUE=19'b0000000_100100111001;
      15'b011_000000100100 : VALUE=19'b0000000_100100111001;
      15'b011_000000100101 : VALUE=19'b0000000_100100111001;
      15'b011_000000100110 : VALUE=19'b0000000_100100111001;
      15'b011_000000100111 : VALUE=19'b0000000_100100111001;
      15'b011_000000101000 : VALUE=19'b0000000_100100111001;
      15'b011_000000101001 : VALUE=19'b0000000_100100111001;
      15'b011_000000101010 : VALUE=19'b0000000_100100111001;
      15'b011_000000101011 : VALUE=19'b0000000_100100111001;
      15'b011_000000101100 : VALUE=19'b0000000_100100111001;
      15'b011_000000101101 : VALUE=19'b0000000_100100111001;
      15'b011_000000101110 : VALUE=19'b0000000_100100111000;
      15'b011_000000101111 : VALUE=19'b0000000_100100111000;
      15'b011_000000110000 : VALUE=19'b0000000_100100111000;
      15'b011_000000110001 : VALUE=19'b0000000_100100111000;
      15'b011_000000110010 : VALUE=19'b0000000_100100111000;
      15'b011_000000110011 : VALUE=19'b0000000_100100111000;
      15'b011_000000110100 : VALUE=19'b0000000_100100111000;
      15'b011_000000110101 : VALUE=19'b0000000_100100111000;
      15'b011_000000110110 : VALUE=19'b0000000_100100111000;
      15'b011_000000110111 : VALUE=19'b0000000_100100111000;
      15'b011_000000111000 : VALUE=19'b0000000_100100110111;
      15'b011_000000111001 : VALUE=19'b0000000_100100110111;
      15'b011_000000111010 : VALUE=19'b0000000_100100110111;
      15'b011_000000111011 : VALUE=19'b0000000_100100110111;
      15'b011_000000111100 : VALUE=19'b0000000_100100110111;
      15'b011_000000111101 : VALUE=19'b0000000_100100110111;
      15'b011_000000111110 : VALUE=19'b0000000_100100110111;
      15'b011_000000111111 : VALUE=19'b0000000_100100110111;
      15'b011_000001000000 : VALUE=19'b0000000_100100110111;
      15'b011_000001000001 : VALUE=19'b0000000_100100110111;
      15'b011_000001000010 : VALUE=19'b0000000_100100110111;
      15'b011_000001000011 : VALUE=19'b0000000_100100110110;
      15'b011_000001000100 : VALUE=19'b0000000_100100110110;
      15'b011_000001000101 : VALUE=19'b0000000_100100110110;
      15'b011_000001000110 : VALUE=19'b0000000_100100110110;
      15'b011_000001000111 : VALUE=19'b0000000_100100110110;
      15'b011_000001001000 : VALUE=19'b0000000_100100110110;
      15'b011_000001001001 : VALUE=19'b0000000_100100110110;
      15'b011_000001001010 : VALUE=19'b0000000_100100110110;
      15'b011_000001001011 : VALUE=19'b0000000_100100110110;
      15'b011_000001001100 : VALUE=19'b0000000_100100110110;
      15'b011_000001001101 : VALUE=19'b0000000_100100110101;
      15'b011_000001001110 : VALUE=19'b0000000_100100110101;
      15'b011_000001001111 : VALUE=19'b0000000_100100110101;
      15'b011_000001010000 : VALUE=19'b0000000_100100110101;
      15'b011_000001010001 : VALUE=19'b0000000_100100110101;
      15'b011_000001010010 : VALUE=19'b0000000_100100110101;
      15'b011_000001010011 : VALUE=19'b0000000_100100110101;
      15'b011_000001010100 : VALUE=19'b0000000_100100110101;
      15'b011_000001010101 : VALUE=19'b0000000_100100110101;
      15'b011_000001010110 : VALUE=19'b0000000_100100110101;
      15'b011_000001010111 : VALUE=19'b0000000_100100110100;
      15'b011_000001011000 : VALUE=19'b0000000_100100110100;
      15'b011_000001011001 : VALUE=19'b0000000_100100110100;
      15'b011_000001011010 : VALUE=19'b0000000_100100110100;
      15'b011_000001011011 : VALUE=19'b0000000_100100110100;
      15'b011_000001011100 : VALUE=19'b0000000_100100110100;
      15'b011_000001011101 : VALUE=19'b0000000_100100110100;
      15'b011_000001011110 : VALUE=19'b0000000_100100110100;
      15'b011_000001011111 : VALUE=19'b0000000_100100110100;
      15'b011_000001100000 : VALUE=19'b0000000_100100110100;
      15'b011_000001100001 : VALUE=19'b0000000_100100110100;
      15'b011_000001100010 : VALUE=19'b0000000_100100110011;
      15'b011_000001100011 : VALUE=19'b0000000_100100110011;
      15'b011_000001100100 : VALUE=19'b0000000_100100110011;
      15'b011_000001100101 : VALUE=19'b0000000_100100110011;
      15'b011_000001100110 : VALUE=19'b0000000_100100110011;
      15'b011_000001100111 : VALUE=19'b0000000_100100110011;
      15'b011_000001101000 : VALUE=19'b0000000_100100110011;
      15'b011_000001101001 : VALUE=19'b0000000_100100110011;
      15'b011_000001101010 : VALUE=19'b0000000_100100110011;
      15'b011_000001101011 : VALUE=19'b0000000_100100110011;
      15'b011_000001101100 : VALUE=19'b0000000_100100110011;
      15'b011_000001101101 : VALUE=19'b0000000_100100110010;
      15'b011_000001101110 : VALUE=19'b0000000_100100110010;
      15'b011_000001101111 : VALUE=19'b0000000_100100110010;
      15'b011_000001110000 : VALUE=19'b0000000_100100110010;
      15'b011_000001110001 : VALUE=19'b0000000_100100110010;
      15'b011_000001110010 : VALUE=19'b0000000_100100110010;
      15'b011_000001110011 : VALUE=19'b0000000_100100110010;
      15'b011_000001110100 : VALUE=19'b0000000_100100110010;
      15'b011_000001110101 : VALUE=19'b0000000_100100110010;
      15'b011_000001110110 : VALUE=19'b0000000_100100110010;
      15'b011_000001110111 : VALUE=19'b0000000_100100110001;
      15'b011_000001111000 : VALUE=19'b0000000_100100110001;
      15'b011_000001111001 : VALUE=19'b0000000_100100110001;
      15'b011_000001111010 : VALUE=19'b0000000_100100110001;
      15'b011_000001111011 : VALUE=19'b0000000_100100110001;
      15'b011_000001111100 : VALUE=19'b0000000_100100110001;
      15'b011_000001111101 : VALUE=19'b0000000_100100110001;
      15'b011_000001111110 : VALUE=19'b0000000_100100110001;
      15'b011_000001111111 : VALUE=19'b0000000_100100110001;
      15'b011_000010000000 : VALUE=19'b0000000_100100110001;
      15'b011_000010000001 : VALUE=19'b0000000_100100110001;
      15'b011_000010000010 : VALUE=19'b0000000_100100110000;
      15'b011_000010000011 : VALUE=19'b0000000_100100110000;
      15'b011_000010000100 : VALUE=19'b0000000_100100110000;
      15'b011_000010000101 : VALUE=19'b0000000_100100110000;
      15'b011_000010000110 : VALUE=19'b0000000_100100110000;
      15'b011_000010000111 : VALUE=19'b0000000_100100110000;
      15'b011_000010001000 : VALUE=19'b0000000_100100110000;
      15'b011_000010001001 : VALUE=19'b0000000_100100110000;
      15'b011_000010001010 : VALUE=19'b0000000_100100110000;
      15'b011_000010001011 : VALUE=19'b0000000_100100110000;
      15'b011_000010001100 : VALUE=19'b0000000_100100101111;
      15'b011_000010001101 : VALUE=19'b0000000_100100101111;
      15'b011_000010001110 : VALUE=19'b0000000_100100101111;
      15'b011_000010001111 : VALUE=19'b0000000_100100101111;
      15'b011_000010010000 : VALUE=19'b0000000_100100101111;
      15'b011_000010010001 : VALUE=19'b0000000_100100101111;
      15'b011_000010010010 : VALUE=19'b0000000_100100101111;
      15'b011_000010010011 : VALUE=19'b0000000_100100101111;
      15'b011_000010010100 : VALUE=19'b0000000_100100101111;
      15'b011_000010010101 : VALUE=19'b0000000_100100101111;
      15'b011_000010010110 : VALUE=19'b0000000_100100101111;
      15'b011_000010010111 : VALUE=19'b0000000_100100101110;
      15'b011_000010011000 : VALUE=19'b0000000_100100101110;
      15'b011_000010011001 : VALUE=19'b0000000_100100101110;
      15'b011_000010011010 : VALUE=19'b0000000_100100101110;
      15'b011_000010011011 : VALUE=19'b0000000_100100101110;
      15'b011_000010011100 : VALUE=19'b0000000_100100101110;
      15'b011_000010011101 : VALUE=19'b0000000_100100101110;
      15'b011_000010011110 : VALUE=19'b0000000_100100101110;
      15'b011_000010011111 : VALUE=19'b0000000_100100101110;
      15'b011_000010100000 : VALUE=19'b0000000_100100101110;
      15'b011_000010100001 : VALUE=19'b0000000_100100101101;
      15'b011_000010100010 : VALUE=19'b0000000_100100101101;
      15'b011_000010100011 : VALUE=19'b0000000_100100101101;
      15'b011_000010100100 : VALUE=19'b0000000_100100101101;
      15'b011_000010100101 : VALUE=19'b0000000_100100101101;
      15'b011_000010100110 : VALUE=19'b0000000_100100101101;
      15'b011_000010100111 : VALUE=19'b0000000_100100101101;
      15'b011_000010101000 : VALUE=19'b0000000_100100101101;
      15'b011_000010101001 : VALUE=19'b0000000_100100101101;
      15'b011_000010101010 : VALUE=19'b0000000_100100101101;
      15'b011_000010101011 : VALUE=19'b0000000_100100101101;
      15'b011_000010101100 : VALUE=19'b0000000_100100101100;
      15'b011_000010101101 : VALUE=19'b0000000_100100101100;
      15'b011_000010101110 : VALUE=19'b0000000_100100101100;
      15'b011_000010101111 : VALUE=19'b0000000_100100101100;
      15'b011_000010110000 : VALUE=19'b0000000_100100101100;
      15'b011_000010110001 : VALUE=19'b0000000_100100101100;
      15'b011_000010110010 : VALUE=19'b0000000_100100101100;
      15'b011_000010110011 : VALUE=19'b0000000_100100101100;
      15'b011_000010110100 : VALUE=19'b0000000_100100101100;
      15'b011_000010110101 : VALUE=19'b0000000_100100101100;
      15'b011_000010110110 : VALUE=19'b0000000_100100101100;
      15'b011_000010110111 : VALUE=19'b0000000_100100101011;
      15'b011_000010111000 : VALUE=19'b0000000_100100101011;
      15'b011_000010111001 : VALUE=19'b0000000_100100101011;
      15'b011_000010111010 : VALUE=19'b0000000_100100101011;
      15'b011_000010111011 : VALUE=19'b0000000_100100101011;
      15'b011_000010111100 : VALUE=19'b0000000_100100101011;
      15'b011_000010111101 : VALUE=19'b0000000_100100101011;
      15'b011_000010111110 : VALUE=19'b0000000_100100101011;
      15'b011_000010111111 : VALUE=19'b0000000_100100101011;
      15'b011_000011000000 : VALUE=19'b0000000_100100101011;
      15'b011_000011000001 : VALUE=19'b0000000_100100101010;
      15'b011_000011000010 : VALUE=19'b0000000_100100101010;
      15'b011_000011000011 : VALUE=19'b0000000_100100101010;
      15'b011_000011000100 : VALUE=19'b0000000_100100101010;
      15'b011_000011000101 : VALUE=19'b0000000_100100101010;
      15'b011_000011000110 : VALUE=19'b0000000_100100101010;
      15'b011_000011000111 : VALUE=19'b0000000_100100101010;
      15'b011_000011001000 : VALUE=19'b0000000_100100101010;
      15'b011_000011001001 : VALUE=19'b0000000_100100101010;
      15'b011_000011001010 : VALUE=19'b0000000_100100101010;
      15'b011_000011001011 : VALUE=19'b0000000_100100101010;
      15'b011_000011001100 : VALUE=19'b0000000_100100101001;
      15'b011_000011001101 : VALUE=19'b0000000_100100101001;
      15'b011_000011001110 : VALUE=19'b0000000_100100101001;
      15'b011_000011001111 : VALUE=19'b0000000_100100101001;
      15'b011_000011010000 : VALUE=19'b0000000_100100101001;
      15'b011_000011010001 : VALUE=19'b0000000_100100101001;
      15'b011_000011010010 : VALUE=19'b0000000_100100101001;
      15'b011_000011010011 : VALUE=19'b0000000_100100101001;
      15'b011_000011010100 : VALUE=19'b0000000_100100101001;
      15'b011_000011010101 : VALUE=19'b0000000_100100101001;
      15'b011_000011010110 : VALUE=19'b0000000_100100101000;
      15'b011_000011010111 : VALUE=19'b0000000_100100101000;
      15'b011_000011011000 : VALUE=19'b0000000_100100101000;
      15'b011_000011011001 : VALUE=19'b0000000_100100101000;
      15'b011_000011011010 : VALUE=19'b0000000_100100101000;
      15'b011_000011011011 : VALUE=19'b0000000_100100101000;
      15'b011_000011011100 : VALUE=19'b0000000_100100101000;
      15'b011_000011011101 : VALUE=19'b0000000_100100101000;
      15'b011_000011011110 : VALUE=19'b0000000_100100101000;
      15'b011_000011011111 : VALUE=19'b0000000_100100101000;
      15'b011_000011100000 : VALUE=19'b0000000_100100101000;
      15'b011_000011100001 : VALUE=19'b0000000_100100100111;
      15'b011_000011100010 : VALUE=19'b0000000_100100100111;
      15'b011_000011100011 : VALUE=19'b0000000_100100100111;
      15'b011_000011100100 : VALUE=19'b0000000_100100100111;
      15'b011_000011100101 : VALUE=19'b0000000_100100100111;
      15'b011_000011100110 : VALUE=19'b0000000_100100100111;
      15'b011_000011100111 : VALUE=19'b0000000_100100100111;
      15'b011_000011101000 : VALUE=19'b0000000_100100100111;
      15'b011_000011101001 : VALUE=19'b0000000_100100100111;
      15'b011_000011101010 : VALUE=19'b0000000_100100100111;
      15'b011_000011101011 : VALUE=19'b0000000_100100100111;
      15'b011_000011101100 : VALUE=19'b0000000_100100100110;
      15'b011_000011101101 : VALUE=19'b0000000_100100100110;
      15'b011_000011101110 : VALUE=19'b0000000_100100100110;
      15'b011_000011101111 : VALUE=19'b0000000_100100100110;
      15'b011_000011110000 : VALUE=19'b0000000_100100100110;
      15'b011_000011110001 : VALUE=19'b0000000_100100100110;
      15'b011_000011110010 : VALUE=19'b0000000_100100100110;
      15'b011_000011110011 : VALUE=19'b0000000_100100100110;
      15'b011_000011110100 : VALUE=19'b0000000_100100100110;
      15'b011_000011110101 : VALUE=19'b0000000_100100100110;
      15'b011_000011110110 : VALUE=19'b0000000_100100100110;
      15'b011_000011110111 : VALUE=19'b0000000_100100100101;
      15'b011_000011111000 : VALUE=19'b0000000_100100100101;
      15'b011_000011111001 : VALUE=19'b0000000_100100100101;
      15'b011_000011111010 : VALUE=19'b0000000_100100100101;
      15'b011_000011111011 : VALUE=19'b0000000_100100100101;
      15'b011_000011111100 : VALUE=19'b0000000_100100100101;
      15'b011_000011111101 : VALUE=19'b0000000_100100100101;
      15'b011_000011111110 : VALUE=19'b0000000_100100100101;
      15'b011_000011111111 : VALUE=19'b0000000_100100100101;
      15'b011_000100000000 : VALUE=19'b0000000_100100100101;
      15'b011_000100000001 : VALUE=19'b0000000_100100100100;
      15'b011_000100000010 : VALUE=19'b0000000_100100100100;
      15'b011_000100000011 : VALUE=19'b0000000_100100100100;
      15'b011_000100000100 : VALUE=19'b0000000_100100100100;
      15'b011_000100000101 : VALUE=19'b0000000_100100100100;
      15'b011_000100000110 : VALUE=19'b0000000_100100100100;
      15'b011_000100000111 : VALUE=19'b0000000_100100100100;
      15'b011_000100001000 : VALUE=19'b0000000_100100100100;
      15'b011_000100001001 : VALUE=19'b0000000_100100100100;
      15'b011_000100001010 : VALUE=19'b0000000_100100100100;
      15'b011_000100001011 : VALUE=19'b0000000_100100100100;
      15'b011_000100001100 : VALUE=19'b0000000_100100100011;
      15'b011_000100001101 : VALUE=19'b0000000_100100100011;
      15'b011_000100001110 : VALUE=19'b0000000_100100100011;
      15'b011_000100001111 : VALUE=19'b0000000_100100100011;
      15'b011_000100010000 : VALUE=19'b0000000_100100100011;
      15'b011_000100010001 : VALUE=19'b0000000_100100100011;
      15'b011_000100010010 : VALUE=19'b0000000_100100100011;
      15'b011_000100010011 : VALUE=19'b0000000_100100100011;
      15'b011_000100010100 : VALUE=19'b0000000_100100100011;
      15'b011_000100010101 : VALUE=19'b0000000_100100100011;
      15'b011_000100010110 : VALUE=19'b0000000_100100100011;
      15'b011_000100010111 : VALUE=19'b0000000_100100100010;
      15'b011_000100011000 : VALUE=19'b0000000_100100100010;
      15'b011_000100011001 : VALUE=19'b0000000_100100100010;
      15'b011_000100011010 : VALUE=19'b0000000_100100100010;
      15'b011_000100011011 : VALUE=19'b0000000_100100100010;
      15'b011_000100011100 : VALUE=19'b0000000_100100100010;
      15'b011_000100011101 : VALUE=19'b0000000_100100100010;
      15'b011_000100011110 : VALUE=19'b0000000_100100100010;
      15'b011_000100011111 : VALUE=19'b0000000_100100100010;
      15'b011_000100100000 : VALUE=19'b0000000_100100100010;
      15'b011_000100100001 : VALUE=19'b0000000_100100100001;
      15'b011_000100100010 : VALUE=19'b0000000_100100100001;
      15'b011_000100100011 : VALUE=19'b0000000_100100100001;
      15'b011_000100100100 : VALUE=19'b0000000_100100100001;
      15'b011_000100100101 : VALUE=19'b0000000_100100100001;
      15'b011_000100100110 : VALUE=19'b0000000_100100100001;
      15'b011_000100100111 : VALUE=19'b0000000_100100100001;
      15'b011_000100101000 : VALUE=19'b0000000_100100100001;
      15'b011_000100101001 : VALUE=19'b0000000_100100100001;
      15'b011_000100101010 : VALUE=19'b0000000_100100100001;
      15'b011_000100101011 : VALUE=19'b0000000_100100100001;
      15'b011_000100101100 : VALUE=19'b0000000_100100100000;
      15'b011_000100101101 : VALUE=19'b0000000_100100100000;
      15'b011_000100101110 : VALUE=19'b0000000_100100100000;
      15'b011_000100101111 : VALUE=19'b0000000_100100100000;
      15'b011_000100110000 : VALUE=19'b0000000_100100100000;
      15'b011_000100110001 : VALUE=19'b0000000_100100100000;
      15'b011_000100110010 : VALUE=19'b0000000_100100100000;
      15'b011_000100110011 : VALUE=19'b0000000_100100100000;
      15'b011_000100110100 : VALUE=19'b0000000_100100100000;
      15'b011_000100110101 : VALUE=19'b0000000_100100100000;
      15'b011_000100110110 : VALUE=19'b0000000_100100100000;
      15'b011_000100110111 : VALUE=19'b0000000_100100011111;
      15'b011_000100111000 : VALUE=19'b0000000_100100011111;
      15'b011_000100111001 : VALUE=19'b0000000_100100011111;
      15'b011_000100111010 : VALUE=19'b0000000_100100011111;
      15'b011_000100111011 : VALUE=19'b0000000_100100011111;
      15'b011_000100111100 : VALUE=19'b0000000_100100011111;
      15'b011_000100111101 : VALUE=19'b0000000_100100011111;
      15'b011_000100111110 : VALUE=19'b0000000_100100011111;
      15'b011_000100111111 : VALUE=19'b0000000_100100011111;
      15'b011_000101000000 : VALUE=19'b0000000_100100011111;
      15'b011_000101000001 : VALUE=19'b0000000_100100011111;
      15'b011_000101000010 : VALUE=19'b0000000_100100011110;
      15'b011_000101000011 : VALUE=19'b0000000_100100011110;
      15'b011_000101000100 : VALUE=19'b0000000_100100011110;
      15'b011_000101000101 : VALUE=19'b0000000_100100011110;
      15'b011_000101000110 : VALUE=19'b0000000_100100011110;
      15'b011_000101000111 : VALUE=19'b0000000_100100011110;
      15'b011_000101001000 : VALUE=19'b0000000_100100011110;
      15'b011_000101001001 : VALUE=19'b0000000_100100011110;
      15'b011_000101001010 : VALUE=19'b0000000_100100011110;
      15'b011_000101001011 : VALUE=19'b0000000_100100011110;
      15'b011_000101001100 : VALUE=19'b0000000_100100011110;
      15'b011_000101001101 : VALUE=19'b0000000_100100011101;
      15'b011_000101001110 : VALUE=19'b0000000_100100011101;
      15'b011_000101001111 : VALUE=19'b0000000_100100011101;
      15'b011_000101010000 : VALUE=19'b0000000_100100011101;
      15'b011_000101010001 : VALUE=19'b0000000_100100011101;
      15'b011_000101010010 : VALUE=19'b0000000_100100011101;
      15'b011_000101010011 : VALUE=19'b0000000_100100011101;
      15'b011_000101010100 : VALUE=19'b0000000_100100011101;
      15'b011_000101010101 : VALUE=19'b0000000_100100011101;
      15'b011_000101010110 : VALUE=19'b0000000_100100011101;
      15'b011_000101010111 : VALUE=19'b0000000_100100011100;
      15'b011_000101011000 : VALUE=19'b0000000_100100011100;
      15'b011_000101011001 : VALUE=19'b0000000_100100011100;
      15'b011_000101011010 : VALUE=19'b0000000_100100011100;
      15'b011_000101011011 : VALUE=19'b0000000_100100011100;
      15'b011_000101011100 : VALUE=19'b0000000_100100011100;
      15'b011_000101011101 : VALUE=19'b0000000_100100011100;
      15'b011_000101011110 : VALUE=19'b0000000_100100011100;
      15'b011_000101011111 : VALUE=19'b0000000_100100011100;
      15'b011_000101100000 : VALUE=19'b0000000_100100011100;
      15'b011_000101100001 : VALUE=19'b0000000_100100011100;
      15'b011_000101100010 : VALUE=19'b0000000_100100011011;
      15'b011_000101100011 : VALUE=19'b0000000_100100011011;
      15'b011_000101100100 : VALUE=19'b0000000_100100011011;
      15'b011_000101100101 : VALUE=19'b0000000_100100011011;
      15'b011_000101100110 : VALUE=19'b0000000_100100011011;
      15'b011_000101100111 : VALUE=19'b0000000_100100011011;
      15'b011_000101101000 : VALUE=19'b0000000_100100011011;
      15'b011_000101101001 : VALUE=19'b0000000_100100011011;
      15'b011_000101101010 : VALUE=19'b0000000_100100011011;
      15'b011_000101101011 : VALUE=19'b0000000_100100011011;
      15'b011_000101101100 : VALUE=19'b0000000_100100011011;
      15'b011_000101101101 : VALUE=19'b0000000_100100011010;
      15'b011_000101101110 : VALUE=19'b0000000_100100011010;
      15'b011_000101101111 : VALUE=19'b0000000_100100011010;
      15'b011_000101110000 : VALUE=19'b0000000_100100011010;
      15'b011_000101110001 : VALUE=19'b0000000_100100011010;
      15'b011_000101110010 : VALUE=19'b0000000_100100011010;
      15'b011_000101110011 : VALUE=19'b0000000_100100011010;
      15'b011_000101110100 : VALUE=19'b0000000_100100011010;
      15'b011_000101110101 : VALUE=19'b0000000_100100011010;
      15'b011_000101110110 : VALUE=19'b0000000_100100011010;
      15'b011_000101110111 : VALUE=19'b0000000_100100011010;
      15'b011_000101111000 : VALUE=19'b0000000_100100011001;
      15'b011_000101111001 : VALUE=19'b0000000_100100011001;
      15'b011_000101111010 : VALUE=19'b0000000_100100011001;
      15'b011_000101111011 : VALUE=19'b0000000_100100011001;
      15'b011_000101111100 : VALUE=19'b0000000_100100011001;
      15'b011_000101111101 : VALUE=19'b0000000_100100011001;
      15'b011_000101111110 : VALUE=19'b0000000_100100011001;
      15'b011_000101111111 : VALUE=19'b0000000_100100011001;
      15'b011_000110000000 : VALUE=19'b0000000_100100011001;
      15'b011_000110000001 : VALUE=19'b0000000_100100011001;
      15'b011_000110000010 : VALUE=19'b0000000_100100011001;
      15'b011_000110000011 : VALUE=19'b0000000_100100011000;
      15'b011_000110000100 : VALUE=19'b0000000_100100011000;
      15'b011_000110000101 : VALUE=19'b0000000_100100011000;
      15'b011_000110000110 : VALUE=19'b0000000_100100011000;
      15'b011_000110000111 : VALUE=19'b0000000_100100011000;
      15'b011_000110001000 : VALUE=19'b0000000_100100011000;
      15'b011_000110001001 : VALUE=19'b0000000_100100011000;
      15'b011_000110001010 : VALUE=19'b0000000_100100011000;
      15'b011_000110001011 : VALUE=19'b0000000_100100011000;
      15'b011_000110001100 : VALUE=19'b0000000_100100011000;
      15'b011_000110001101 : VALUE=19'b0000000_100100011000;
      15'b011_000110001110 : VALUE=19'b0000000_100100010111;
      15'b011_000110001111 : VALUE=19'b0000000_100100010111;
      15'b011_000110010000 : VALUE=19'b0000000_100100010111;
      15'b011_000110010001 : VALUE=19'b0000000_100100010111;
      15'b011_000110010010 : VALUE=19'b0000000_100100010111;
      15'b011_000110010011 : VALUE=19'b0000000_100100010111;
      15'b011_000110010100 : VALUE=19'b0000000_100100010111;
      15'b011_000110010101 : VALUE=19'b0000000_100100010111;
      15'b011_000110010110 : VALUE=19'b0000000_100100010111;
      15'b011_000110010111 : VALUE=19'b0000000_100100010111;
      15'b011_000110011000 : VALUE=19'b0000000_100100010111;
      15'b011_000110011001 : VALUE=19'b0000000_100100010110;
      15'b011_000110011010 : VALUE=19'b0000000_100100010110;
      15'b011_000110011011 : VALUE=19'b0000000_100100010110;
      15'b011_000110011100 : VALUE=19'b0000000_100100010110;
      15'b011_000110011101 : VALUE=19'b0000000_100100010110;
      15'b011_000110011110 : VALUE=19'b0000000_100100010110;
      15'b011_000110011111 : VALUE=19'b0000000_100100010110;
      15'b011_000110100000 : VALUE=19'b0000000_100100010110;
      15'b011_000110100001 : VALUE=19'b0000000_100100010110;
      15'b011_000110100010 : VALUE=19'b0000000_100100010110;
      15'b011_000110100011 : VALUE=19'b0000000_100100010110;
      15'b011_000110100100 : VALUE=19'b0000000_100100010101;
      15'b011_000110100101 : VALUE=19'b0000000_100100010101;
      15'b011_000110100110 : VALUE=19'b0000000_100100010101;
      15'b011_000110100111 : VALUE=19'b0000000_100100010101;
      15'b011_000110101000 : VALUE=19'b0000000_100100010101;
      15'b011_000110101001 : VALUE=19'b0000000_100100010101;
      15'b011_000110101010 : VALUE=19'b0000000_100100010101;
      15'b011_000110101011 : VALUE=19'b0000000_100100010101;
      15'b011_000110101100 : VALUE=19'b0000000_100100010101;
      15'b011_000110101101 : VALUE=19'b0000000_100100010101;
      15'b011_000110101110 : VALUE=19'b0000000_100100010101;
      15'b011_000110101111 : VALUE=19'b0000000_100100010100;
      15'b011_000110110000 : VALUE=19'b0000000_100100010100;
      15'b011_000110110001 : VALUE=19'b0000000_100100010100;
      15'b011_000110110010 : VALUE=19'b0000000_100100010100;
      15'b011_000110110011 : VALUE=19'b0000000_100100010100;
      15'b011_000110110100 : VALUE=19'b0000000_100100010100;
      15'b011_000110110101 : VALUE=19'b0000000_100100010100;
      15'b011_000110110110 : VALUE=19'b0000000_100100010100;
      15'b011_000110110111 : VALUE=19'b0000000_100100010100;
      15'b011_000110111000 : VALUE=19'b0000000_100100010100;
      15'b011_000110111001 : VALUE=19'b0000000_100100010100;
      15'b011_000110111010 : VALUE=19'b0000000_100100010011;
      15'b011_000110111011 : VALUE=19'b0000000_100100010011;
      15'b011_000110111100 : VALUE=19'b0000000_100100010011;
      15'b011_000110111101 : VALUE=19'b0000000_100100010011;
      15'b011_000110111110 : VALUE=19'b0000000_100100010011;
      15'b011_000110111111 : VALUE=19'b0000000_100100010011;
      15'b011_000111000000 : VALUE=19'b0000000_100100010011;
      15'b011_000111000001 : VALUE=19'b0000000_100100010011;
      15'b011_000111000010 : VALUE=19'b0000000_100100010011;
      15'b011_000111000011 : VALUE=19'b0000000_100100010011;
      15'b011_000111000100 : VALUE=19'b0000000_100100010010;
      15'b011_000111000101 : VALUE=19'b0000000_100100010010;
      15'b011_000111000110 : VALUE=19'b0000000_100100010010;
      15'b011_000111000111 : VALUE=19'b0000000_100100010010;
      15'b011_000111001000 : VALUE=19'b0000000_100100010010;
      15'b011_000111001001 : VALUE=19'b0000000_100100010010;
      15'b011_000111001010 : VALUE=19'b0000000_100100010010;
      15'b011_000111001011 : VALUE=19'b0000000_100100010010;
      15'b011_000111001100 : VALUE=19'b0000000_100100010010;
      15'b011_000111001101 : VALUE=19'b0000000_100100010010;
      15'b011_000111001110 : VALUE=19'b0000000_100100010010;
      15'b011_000111001111 : VALUE=19'b0000000_100100010001;
      15'b011_000111010000 : VALUE=19'b0000000_100100010001;
      15'b011_000111010001 : VALUE=19'b0000000_100100010001;
      15'b011_000111010010 : VALUE=19'b0000000_100100010001;
      15'b011_000111010011 : VALUE=19'b0000000_100100010001;
      15'b011_000111010100 : VALUE=19'b0000000_100100010001;
      15'b011_000111010101 : VALUE=19'b0000000_100100010001;
      15'b011_000111010110 : VALUE=19'b0000000_100100010001;
      15'b011_000111010111 : VALUE=19'b0000000_100100010001;
      15'b011_000111011000 : VALUE=19'b0000000_100100010001;
      15'b011_000111011001 : VALUE=19'b0000000_100100010001;
      15'b011_000111011010 : VALUE=19'b0000000_100100010000;
      15'b011_000111011011 : VALUE=19'b0000000_100100010000;
      15'b011_000111011100 : VALUE=19'b0000000_100100010000;
      15'b011_000111011101 : VALUE=19'b0000000_100100010000;
      15'b011_000111011110 : VALUE=19'b0000000_100100010000;
      15'b011_000111011111 : VALUE=19'b0000000_100100010000;
      15'b011_000111100000 : VALUE=19'b0000000_100100010000;
      15'b011_000111100001 : VALUE=19'b0000000_100100010000;
      15'b011_000111100010 : VALUE=19'b0000000_100100010000;
      15'b011_000111100011 : VALUE=19'b0000000_100100010000;
      15'b011_000111100100 : VALUE=19'b0000000_100100010000;
      15'b011_000111100101 : VALUE=19'b0000000_100100001111;
      15'b011_000111100110 : VALUE=19'b0000000_100100001111;
      15'b011_000111100111 : VALUE=19'b0000000_100100001111;
      15'b011_000111101000 : VALUE=19'b0000000_100100001111;
      15'b011_000111101001 : VALUE=19'b0000000_100100001111;
      15'b011_000111101010 : VALUE=19'b0000000_100100001111;
      15'b011_000111101011 : VALUE=19'b0000000_100100001111;
      15'b011_000111101100 : VALUE=19'b0000000_100100001111;
      15'b011_000111101101 : VALUE=19'b0000000_100100001111;
      15'b011_000111101110 : VALUE=19'b0000000_100100001111;
      15'b011_000111101111 : VALUE=19'b0000000_100100001111;
      15'b011_000111110000 : VALUE=19'b0000000_100100001110;
      15'b011_000111110001 : VALUE=19'b0000000_100100001110;
      15'b011_000111110010 : VALUE=19'b0000000_100100001110;
      15'b011_000111110011 : VALUE=19'b0000000_100100001110;
      15'b011_000111110100 : VALUE=19'b0000000_100100001110;
      15'b011_000111110101 : VALUE=19'b0000000_100100001110;
      15'b011_000111110110 : VALUE=19'b0000000_100100001110;
      15'b011_000111110111 : VALUE=19'b0000000_100100001110;
      15'b011_000111111000 : VALUE=19'b0000000_100100001110;
      15'b011_000111111001 : VALUE=19'b0000000_100100001110;
      15'b011_000111111010 : VALUE=19'b0000000_100100001110;
      15'b011_000111111011 : VALUE=19'b0000000_100100001110;
      15'b011_000111111100 : VALUE=19'b0000000_100100001101;
      15'b011_000111111101 : VALUE=19'b0000000_100100001101;
      15'b011_000111111110 : VALUE=19'b0000000_100100001101;
      15'b011_000111111111 : VALUE=19'b0000000_100100001101;
      15'b011_001000000000 : VALUE=19'b0000000_100100001101;
      15'b011_001000000001 : VALUE=19'b0000000_100100001101;
      15'b011_001000000010 : VALUE=19'b0000000_100100001101;
      15'b011_001000000011 : VALUE=19'b0000000_100100001101;
      15'b011_001000000100 : VALUE=19'b0000000_100100001101;
      15'b011_001000000101 : VALUE=19'b0000000_100100001101;
      15'b011_001000000110 : VALUE=19'b0000000_100100001101;
      15'b011_001000000111 : VALUE=19'b0000000_100100001100;
      15'b011_001000001000 : VALUE=19'b0000000_100100001100;
      15'b011_001000001001 : VALUE=19'b0000000_100100001100;
      15'b011_001000001010 : VALUE=19'b0000000_100100001100;
      15'b011_001000001011 : VALUE=19'b0000000_100100001100;
      15'b011_001000001100 : VALUE=19'b0000000_100100001100;
      15'b011_001000001101 : VALUE=19'b0000000_100100001100;
      15'b011_001000001110 : VALUE=19'b0000000_100100001100;
      15'b011_001000001111 : VALUE=19'b0000000_100100001100;
      15'b011_001000010000 : VALUE=19'b0000000_100100001100;
      15'b011_001000010001 : VALUE=19'b0000000_100100001100;
      15'b011_001000010010 : VALUE=19'b0000000_100100001011;
      15'b011_001000010011 : VALUE=19'b0000000_100100001011;
      15'b011_001000010100 : VALUE=19'b0000000_100100001011;
      15'b011_001000010101 : VALUE=19'b0000000_100100001011;
      15'b011_001000010110 : VALUE=19'b0000000_100100001011;
      15'b011_001000010111 : VALUE=19'b0000000_100100001011;
      15'b011_001000011000 : VALUE=19'b0000000_100100001011;
      15'b011_001000011001 : VALUE=19'b0000000_100100001011;
      15'b011_001000011010 : VALUE=19'b0000000_100100001011;
      15'b011_001000011011 : VALUE=19'b0000000_100100001011;
      15'b011_001000011100 : VALUE=19'b0000000_100100001011;
      15'b011_001000011101 : VALUE=19'b0000000_100100001010;
      15'b011_001000011110 : VALUE=19'b0000000_100100001010;
      15'b011_001000011111 : VALUE=19'b0000000_100100001010;
      15'b011_001000100000 : VALUE=19'b0000000_100100001010;
      15'b011_001000100001 : VALUE=19'b0000000_100100001010;
      15'b011_001000100010 : VALUE=19'b0000000_100100001010;
      15'b011_001000100011 : VALUE=19'b0000000_100100001010;
      15'b011_001000100100 : VALUE=19'b0000000_100100001010;
      15'b011_001000100101 : VALUE=19'b0000000_100100001010;
      15'b011_001000100110 : VALUE=19'b0000000_100100001010;
      15'b011_001000100111 : VALUE=19'b0000000_100100001010;
      15'b011_001000101000 : VALUE=19'b0000000_100100001001;
      15'b011_001000101001 : VALUE=19'b0000000_100100001001;
      15'b011_001000101010 : VALUE=19'b0000000_100100001001;
      15'b011_001000101011 : VALUE=19'b0000000_100100001001;
      15'b011_001000101100 : VALUE=19'b0000000_100100001001;
      15'b011_001000101101 : VALUE=19'b0000000_100100001001;
      15'b011_001000101110 : VALUE=19'b0000000_100100001001;
      15'b011_001000101111 : VALUE=19'b0000000_100100001001;
      15'b011_001000110000 : VALUE=19'b0000000_100100001001;
      15'b011_001000110001 : VALUE=19'b0000000_100100001001;
      15'b011_001000110010 : VALUE=19'b0000000_100100001001;
      15'b011_001000110011 : VALUE=19'b0000000_100100001000;
      15'b011_001000110100 : VALUE=19'b0000000_100100001000;
      15'b011_001000110101 : VALUE=19'b0000000_100100001000;
      15'b011_001000110110 : VALUE=19'b0000000_100100001000;
      15'b011_001000110111 : VALUE=19'b0000000_100100001000;
      15'b011_001000111000 : VALUE=19'b0000000_100100001000;
      15'b011_001000111001 : VALUE=19'b0000000_100100001000;
      15'b011_001000111010 : VALUE=19'b0000000_100100001000;
      15'b011_001000111011 : VALUE=19'b0000000_100100001000;
      15'b011_001000111100 : VALUE=19'b0000000_100100001000;
      15'b011_001000111101 : VALUE=19'b0000000_100100001000;
      15'b011_001000111110 : VALUE=19'b0000000_100100000111;
      15'b011_001000111111 : VALUE=19'b0000000_100100000111;
      15'b011_001001000000 : VALUE=19'b0000000_100100000111;
      15'b011_001001000001 : VALUE=19'b0000000_100100000111;
      15'b011_001001000010 : VALUE=19'b0000000_100100000111;
      15'b011_001001000011 : VALUE=19'b0000000_100100000111;
      15'b011_001001000100 : VALUE=19'b0000000_100100000111;
      15'b011_001001000101 : VALUE=19'b0000000_100100000111;
      15'b011_001001000110 : VALUE=19'b0000000_100100000111;
      15'b011_001001000111 : VALUE=19'b0000000_100100000111;
      15'b011_001001001000 : VALUE=19'b0000000_100100000111;
      15'b011_001001001001 : VALUE=19'b0000000_100100000110;
      15'b011_001001001010 : VALUE=19'b0000000_100100000110;
      15'b011_001001001011 : VALUE=19'b0000000_100100000110;
      15'b011_001001001100 : VALUE=19'b0000000_100100000110;
      15'b011_001001001101 : VALUE=19'b0000000_100100000110;
      15'b011_001001001110 : VALUE=19'b0000000_100100000110;
      15'b011_001001001111 : VALUE=19'b0000000_100100000110;
      15'b011_001001010000 : VALUE=19'b0000000_100100000110;
      15'b011_001001010001 : VALUE=19'b0000000_100100000110;
      15'b011_001001010010 : VALUE=19'b0000000_100100000110;
      15'b011_001001010011 : VALUE=19'b0000000_100100000110;
      15'b011_001001010100 : VALUE=19'b0000000_100100000101;
      15'b011_001001010101 : VALUE=19'b0000000_100100000101;
      15'b011_001001010110 : VALUE=19'b0000000_100100000101;
      15'b011_001001010111 : VALUE=19'b0000000_100100000101;
      15'b011_001001011000 : VALUE=19'b0000000_100100000101;
      15'b011_001001011001 : VALUE=19'b0000000_100100000101;
      15'b011_001001011010 : VALUE=19'b0000000_100100000101;
      15'b011_001001011011 : VALUE=19'b0000000_100100000101;
      15'b011_001001011100 : VALUE=19'b0000000_100100000101;
      15'b011_001001011101 : VALUE=19'b0000000_100100000101;
      15'b011_001001011110 : VALUE=19'b0000000_100100000101;
      15'b011_001001011111 : VALUE=19'b0000000_100100000100;
      15'b011_001001100000 : VALUE=19'b0000000_100100000100;
      15'b011_001001100001 : VALUE=19'b0000000_100100000100;
      15'b011_001001100010 : VALUE=19'b0000000_100100000100;
      15'b011_001001100011 : VALUE=19'b0000000_100100000100;
      15'b011_001001100100 : VALUE=19'b0000000_100100000100;
      15'b011_001001100101 : VALUE=19'b0000000_100100000100;
      15'b011_001001100110 : VALUE=19'b0000000_100100000100;
      15'b011_001001100111 : VALUE=19'b0000000_100100000100;
      15'b011_001001101000 : VALUE=19'b0000000_100100000100;
      15'b011_001001101001 : VALUE=19'b0000000_100100000100;
      15'b011_001001101010 : VALUE=19'b0000000_100100000100;
      15'b011_001001101011 : VALUE=19'b0000000_100100000011;
      15'b011_001001101100 : VALUE=19'b0000000_100100000011;
      15'b011_001001101101 : VALUE=19'b0000000_100100000011;
      15'b011_001001101110 : VALUE=19'b0000000_100100000011;
      15'b011_001001101111 : VALUE=19'b0000000_100100000011;
      15'b011_001001110000 : VALUE=19'b0000000_100100000011;
      15'b011_001001110001 : VALUE=19'b0000000_100100000011;
      15'b011_001001110010 : VALUE=19'b0000000_100100000011;
      15'b011_001001110011 : VALUE=19'b0000000_100100000011;
      15'b011_001001110100 : VALUE=19'b0000000_100100000011;
      15'b011_001001110101 : VALUE=19'b0000000_100100000011;
      15'b011_001001110110 : VALUE=19'b0000000_100100000010;
      15'b011_001001110111 : VALUE=19'b0000000_100100000010;
      15'b011_001001111000 : VALUE=19'b0000000_100100000010;
      15'b011_001001111001 : VALUE=19'b0000000_100100000010;
      15'b011_001001111010 : VALUE=19'b0000000_100100000010;
      15'b011_001001111011 : VALUE=19'b0000000_100100000010;
      15'b011_001001111100 : VALUE=19'b0000000_100100000010;
      15'b011_001001111101 : VALUE=19'b0000000_100100000010;
      15'b011_001001111110 : VALUE=19'b0000000_100100000010;
      15'b011_001001111111 : VALUE=19'b0000000_100100000010;
      15'b011_001010000000 : VALUE=19'b0000000_100100000010;
      15'b011_001010000001 : VALUE=19'b0000000_100100000001;
      15'b011_001010000010 : VALUE=19'b0000000_100100000001;
      15'b011_001010000011 : VALUE=19'b0000000_100100000001;
      15'b011_001010000100 : VALUE=19'b0000000_100100000001;
      15'b011_001010000101 : VALUE=19'b0000000_100100000001;
      15'b011_001010000110 : VALUE=19'b0000000_100100000001;
      15'b011_001010000111 : VALUE=19'b0000000_100100000001;
      15'b011_001010001000 : VALUE=19'b0000000_100100000001;
      15'b011_001010001001 : VALUE=19'b0000000_100100000001;
      15'b011_001010001010 : VALUE=19'b0000000_100100000001;
      15'b011_001010001011 : VALUE=19'b0000000_100100000001;
      15'b011_001010001100 : VALUE=19'b0000000_100100000000;
      15'b011_001010001101 : VALUE=19'b0000000_100100000000;
      15'b011_001010001110 : VALUE=19'b0000000_100100000000;
      15'b011_001010001111 : VALUE=19'b0000000_100100000000;
      15'b011_001010010000 : VALUE=19'b0000000_100100000000;
      15'b011_001010010001 : VALUE=19'b0000000_100100000000;
      15'b011_001010010010 : VALUE=19'b0000000_100100000000;
      15'b011_001010010011 : VALUE=19'b0000000_100100000000;
      15'b011_001010010100 : VALUE=19'b0000000_100100000000;
      15'b011_001010010101 : VALUE=19'b0000000_100100000000;
      15'b011_001010010110 : VALUE=19'b0000000_100100000000;
      15'b011_001010010111 : VALUE=19'b0000000_100100000000;
      15'b011_001010011000 : VALUE=19'b0000000_100011111111;
      15'b011_001010011001 : VALUE=19'b0000000_100011111111;
      15'b011_001010011010 : VALUE=19'b0000000_100011111111;
      15'b011_001010011011 : VALUE=19'b0000000_100011111111;
      15'b011_001010011100 : VALUE=19'b0000000_100011111111;
      15'b011_001010011101 : VALUE=19'b0000000_100011111111;
      15'b011_001010011110 : VALUE=19'b0000000_100011111111;
      15'b011_001010011111 : VALUE=19'b0000000_100011111111;
      15'b011_001010100000 : VALUE=19'b0000000_100011111111;
      15'b011_001010100001 : VALUE=19'b0000000_100011111111;
      15'b011_001010100010 : VALUE=19'b0000000_100011111111;
      15'b011_001010100011 : VALUE=19'b0000000_100011111110;
      15'b011_001010100100 : VALUE=19'b0000000_100011111110;
      15'b011_001010100101 : VALUE=19'b0000000_100011111110;
      15'b011_001010100110 : VALUE=19'b0000000_100011111110;
      15'b011_001010100111 : VALUE=19'b0000000_100011111110;
      15'b011_001010101000 : VALUE=19'b0000000_100011111110;
      15'b011_001010101001 : VALUE=19'b0000000_100011111110;
      15'b011_001010101010 : VALUE=19'b0000000_100011111110;
      15'b011_001010101011 : VALUE=19'b0000000_100011111110;
      15'b011_001010101100 : VALUE=19'b0000000_100011111110;
      15'b011_001010101101 : VALUE=19'b0000000_100011111110;
      15'b011_001010101110 : VALUE=19'b0000000_100011111101;
      15'b011_001010101111 : VALUE=19'b0000000_100011111101;
      15'b011_001010110000 : VALUE=19'b0000000_100011111101;
      15'b011_001010110001 : VALUE=19'b0000000_100011111101;
      15'b011_001010110010 : VALUE=19'b0000000_100011111101;
      15'b011_001010110011 : VALUE=19'b0000000_100011111101;
      15'b011_001010110100 : VALUE=19'b0000000_100011111101;
      15'b011_001010110101 : VALUE=19'b0000000_100011111101;
      15'b011_001010110110 : VALUE=19'b0000000_100011111101;
      15'b011_001010110111 : VALUE=19'b0000000_100011111101;
      15'b011_001010111000 : VALUE=19'b0000000_100011111101;
      15'b011_001010111001 : VALUE=19'b0000000_100011111100;
      15'b011_001010111010 : VALUE=19'b0000000_100011111100;
      15'b011_001010111011 : VALUE=19'b0000000_100011111100;
      15'b011_001010111100 : VALUE=19'b0000000_100011111100;
      15'b011_001010111101 : VALUE=19'b0000000_100011111100;
      15'b011_001010111110 : VALUE=19'b0000000_100011111100;
      15'b011_001010111111 : VALUE=19'b0000000_100011111100;
      15'b011_001011000000 : VALUE=19'b0000000_100011111100;
      15'b011_001011000001 : VALUE=19'b0000000_100011111100;
      15'b011_001011000010 : VALUE=19'b0000000_100011111100;
      15'b011_001011000011 : VALUE=19'b0000000_100011111100;
      15'b011_001011000100 : VALUE=19'b0000000_100011111100;
      15'b011_001011000101 : VALUE=19'b0000000_100011111011;
      15'b011_001011000110 : VALUE=19'b0000000_100011111011;
      15'b011_001011000111 : VALUE=19'b0000000_100011111011;
      15'b011_001011001000 : VALUE=19'b0000000_100011111011;
      15'b011_001011001001 : VALUE=19'b0000000_100011111011;
      15'b011_001011001010 : VALUE=19'b0000000_100011111011;
      15'b011_001011001011 : VALUE=19'b0000000_100011111011;
      15'b011_001011001100 : VALUE=19'b0000000_100011111011;
      15'b011_001011001101 : VALUE=19'b0000000_100011111011;
      15'b011_001011001110 : VALUE=19'b0000000_100011111011;
      15'b011_001011001111 : VALUE=19'b0000000_100011111011;
      15'b011_001011010000 : VALUE=19'b0000000_100011111010;
      15'b011_001011010001 : VALUE=19'b0000000_100011111010;
      15'b011_001011010010 : VALUE=19'b0000000_100011111010;
      15'b011_001011010011 : VALUE=19'b0000000_100011111010;
      15'b011_001011010100 : VALUE=19'b0000000_100011111010;
      15'b011_001011010101 : VALUE=19'b0000000_100011111010;
      15'b011_001011010110 : VALUE=19'b0000000_100011111010;
      15'b011_001011010111 : VALUE=19'b0000000_100011111010;
      15'b011_001011011000 : VALUE=19'b0000000_100011111010;
      15'b011_001011011001 : VALUE=19'b0000000_100011111010;
      15'b011_001011011010 : VALUE=19'b0000000_100011111010;
      15'b011_001011011011 : VALUE=19'b0000000_100011111001;
      15'b011_001011011100 : VALUE=19'b0000000_100011111001;
      15'b011_001011011101 : VALUE=19'b0000000_100011111001;
      15'b011_001011011110 : VALUE=19'b0000000_100011111001;
      15'b011_001011011111 : VALUE=19'b0000000_100011111001;
      15'b011_001011100000 : VALUE=19'b0000000_100011111001;
      15'b011_001011100001 : VALUE=19'b0000000_100011111001;
      15'b011_001011100010 : VALUE=19'b0000000_100011111001;
      15'b011_001011100011 : VALUE=19'b0000000_100011111001;
      15'b011_001011100100 : VALUE=19'b0000000_100011111001;
      15'b011_001011100101 : VALUE=19'b0000000_100011111001;
      15'b011_001011100110 : VALUE=19'b0000000_100011111001;
      15'b011_001011100111 : VALUE=19'b0000000_100011111000;
      15'b011_001011101000 : VALUE=19'b0000000_100011111000;
      15'b011_001011101001 : VALUE=19'b0000000_100011111000;
      15'b011_001011101010 : VALUE=19'b0000000_100011111000;
      15'b011_001011101011 : VALUE=19'b0000000_100011111000;
      15'b011_001011101100 : VALUE=19'b0000000_100011111000;
      15'b011_001011101101 : VALUE=19'b0000000_100011111000;
      15'b011_001011101110 : VALUE=19'b0000000_100011111000;
      15'b011_001011101111 : VALUE=19'b0000000_100011111000;
      15'b011_001011110000 : VALUE=19'b0000000_100011111000;
      15'b011_001011110001 : VALUE=19'b0000000_100011111000;
      15'b011_001011110010 : VALUE=19'b0000000_100011110111;
      15'b011_001011110011 : VALUE=19'b0000000_100011110111;
      15'b011_001011110100 : VALUE=19'b0000000_100011110111;
      15'b011_001011110101 : VALUE=19'b0000000_100011110111;
      15'b011_001011110110 : VALUE=19'b0000000_100011110111;
      15'b011_001011110111 : VALUE=19'b0000000_100011110111;
      15'b011_001011111000 : VALUE=19'b0000000_100011110111;
      15'b011_001011111001 : VALUE=19'b0000000_100011110111;
      15'b011_001011111010 : VALUE=19'b0000000_100011110111;
      15'b011_001011111011 : VALUE=19'b0000000_100011110111;
      15'b011_001011111100 : VALUE=19'b0000000_100011110111;
      15'b011_001011111101 : VALUE=19'b0000000_100011110110;
      15'b011_001011111110 : VALUE=19'b0000000_100011110110;
      15'b011_001011111111 : VALUE=19'b0000000_100011110110;
      15'b011_001100000000 : VALUE=19'b0000000_100011110110;
      15'b011_001100000001 : VALUE=19'b0000000_100011110110;
      15'b011_001100000010 : VALUE=19'b0000000_100011110110;
      15'b011_001100000011 : VALUE=19'b0000000_100011110110;
      15'b011_001100000100 : VALUE=19'b0000000_100011110110;
      15'b011_001100000101 : VALUE=19'b0000000_100011110110;
      15'b011_001100000110 : VALUE=19'b0000000_100011110110;
      15'b011_001100000111 : VALUE=19'b0000000_100011110110;
      15'b011_001100001000 : VALUE=19'b0000000_100011110110;
      15'b011_001100001001 : VALUE=19'b0000000_100011110101;
      15'b011_001100001010 : VALUE=19'b0000000_100011110101;
      15'b011_001100001011 : VALUE=19'b0000000_100011110101;
      15'b011_001100001100 : VALUE=19'b0000000_100011110101;
      15'b011_001100001101 : VALUE=19'b0000000_100011110101;
      15'b011_001100001110 : VALUE=19'b0000000_100011110101;
      15'b011_001100001111 : VALUE=19'b0000000_100011110101;
      15'b011_001100010000 : VALUE=19'b0000000_100011110101;
      15'b011_001100010001 : VALUE=19'b0000000_100011110101;
      15'b011_001100010010 : VALUE=19'b0000000_100011110101;
      15'b011_001100010011 : VALUE=19'b0000000_100011110101;
      15'b011_001100010100 : VALUE=19'b0000000_100011110100;
      15'b011_001100010101 : VALUE=19'b0000000_100011110100;
      15'b011_001100010110 : VALUE=19'b0000000_100011110100;
      15'b011_001100010111 : VALUE=19'b0000000_100011110100;
      15'b011_001100011000 : VALUE=19'b0000000_100011110100;
      15'b011_001100011001 : VALUE=19'b0000000_100011110100;
      15'b011_001100011010 : VALUE=19'b0000000_100011110100;
      15'b011_001100011011 : VALUE=19'b0000000_100011110100;
      15'b011_001100011100 : VALUE=19'b0000000_100011110100;
      15'b011_001100011101 : VALUE=19'b0000000_100011110100;
      15'b011_001100011110 : VALUE=19'b0000000_100011110100;
      15'b011_001100011111 : VALUE=19'b0000000_100011110100;
      15'b011_001100100000 : VALUE=19'b0000000_100011110011;
      15'b011_001100100001 : VALUE=19'b0000000_100011110011;
      15'b011_001100100010 : VALUE=19'b0000000_100011110011;
      15'b011_001100100011 : VALUE=19'b0000000_100011110011;
      15'b011_001100100100 : VALUE=19'b0000000_100011110011;
      15'b011_001100100101 : VALUE=19'b0000000_100011110011;
      15'b011_001100100110 : VALUE=19'b0000000_100011110011;
      15'b011_001100100111 : VALUE=19'b0000000_100011110011;
      15'b011_001100101000 : VALUE=19'b0000000_100011110011;
      15'b011_001100101001 : VALUE=19'b0000000_100011110011;
      15'b011_001100101010 : VALUE=19'b0000000_100011110011;
      15'b011_001100101011 : VALUE=19'b0000000_100011110010;
      15'b011_001100101100 : VALUE=19'b0000000_100011110010;
      15'b011_001100101101 : VALUE=19'b0000000_100011110010;
      15'b011_001100101110 : VALUE=19'b0000000_100011110010;
      15'b011_001100101111 : VALUE=19'b0000000_100011110010;
      15'b011_001100110000 : VALUE=19'b0000000_100011110010;
      15'b011_001100110001 : VALUE=19'b0000000_100011110010;
      15'b011_001100110010 : VALUE=19'b0000000_100011110010;
      15'b011_001100110011 : VALUE=19'b0000000_100011110010;
      15'b011_001100110100 : VALUE=19'b0000000_100011110010;
      15'b011_001100110101 : VALUE=19'b0000000_100011110010;
      15'b011_001100110110 : VALUE=19'b0000000_100011110001;
      15'b011_001100110111 : VALUE=19'b0000000_100011110001;
      15'b011_001100111000 : VALUE=19'b0000000_100011110001;
      15'b011_001100111001 : VALUE=19'b0000000_100011110001;
      15'b011_001100111010 : VALUE=19'b0000000_100011110001;
      15'b011_001100111011 : VALUE=19'b0000000_100011110001;
      15'b011_001100111100 : VALUE=19'b0000000_100011110001;
      15'b011_001100111101 : VALUE=19'b0000000_100011110001;
      15'b011_001100111110 : VALUE=19'b0000000_100011110001;
      15'b011_001100111111 : VALUE=19'b0000000_100011110001;
      15'b011_001101000000 : VALUE=19'b0000000_100011110001;
      15'b011_001101000001 : VALUE=19'b0000000_100011110001;
      15'b011_001101000010 : VALUE=19'b0000000_100011110000;
      15'b011_001101000011 : VALUE=19'b0000000_100011110000;
      15'b011_001101000100 : VALUE=19'b0000000_100011110000;
      15'b011_001101000101 : VALUE=19'b0000000_100011110000;
      15'b011_001101000110 : VALUE=19'b0000000_100011110000;
      15'b011_001101000111 : VALUE=19'b0000000_100011110000;
      15'b011_001101001000 : VALUE=19'b0000000_100011110000;
      15'b011_001101001001 : VALUE=19'b0000000_100011110000;
      15'b011_001101001010 : VALUE=19'b0000000_100011110000;
      15'b011_001101001011 : VALUE=19'b0000000_100011110000;
      15'b011_001101001100 : VALUE=19'b0000000_100011110000;
      15'b011_001101001101 : VALUE=19'b0000000_100011101111;
      15'b011_001101001110 : VALUE=19'b0000000_100011101111;
      15'b011_001101001111 : VALUE=19'b0000000_100011101111;
      15'b011_001101010000 : VALUE=19'b0000000_100011101111;
      15'b011_001101010001 : VALUE=19'b0000000_100011101111;
      15'b011_001101010010 : VALUE=19'b0000000_100011101111;
      15'b011_001101010011 : VALUE=19'b0000000_100011101111;
      15'b011_001101010100 : VALUE=19'b0000000_100011101111;
      15'b011_001101010101 : VALUE=19'b0000000_100011101111;
      15'b011_001101010110 : VALUE=19'b0000000_100011101111;
      15'b011_001101010111 : VALUE=19'b0000000_100011101111;
      15'b011_001101011000 : VALUE=19'b0000000_100011101111;
      15'b011_001101011001 : VALUE=19'b0000000_100011101110;
      15'b011_001101011010 : VALUE=19'b0000000_100011101110;
      15'b011_001101011011 : VALUE=19'b0000000_100011101110;
      15'b011_001101011100 : VALUE=19'b0000000_100011101110;
      15'b011_001101011101 : VALUE=19'b0000000_100011101110;
      15'b011_001101011110 : VALUE=19'b0000000_100011101110;
      15'b011_001101011111 : VALUE=19'b0000000_100011101110;
      15'b011_001101100000 : VALUE=19'b0000000_100011101110;
      15'b011_001101100001 : VALUE=19'b0000000_100011101110;
      15'b011_001101100010 : VALUE=19'b0000000_100011101110;
      15'b011_001101100011 : VALUE=19'b0000000_100011101110;
      15'b011_001101100100 : VALUE=19'b0000000_100011101101;
      15'b011_001101100101 : VALUE=19'b0000000_100011101101;
      15'b011_001101100110 : VALUE=19'b0000000_100011101101;
      15'b011_001101100111 : VALUE=19'b0000000_100011101101;
      15'b011_001101101000 : VALUE=19'b0000000_100011101101;
      15'b011_001101101001 : VALUE=19'b0000000_100011101101;
      15'b011_001101101010 : VALUE=19'b0000000_100011101101;
      15'b011_001101101011 : VALUE=19'b0000000_100011101101;
      15'b011_001101101100 : VALUE=19'b0000000_100011101101;
      15'b011_001101101101 : VALUE=19'b0000000_100011101101;
      15'b011_001101101110 : VALUE=19'b0000000_100011101101;
      15'b011_001101101111 : VALUE=19'b0000000_100011101101;
      15'b011_001101110000 : VALUE=19'b0000000_100011101100;
      15'b011_001101110001 : VALUE=19'b0000000_100011101100;
      15'b011_001101110010 : VALUE=19'b0000000_100011101100;
      15'b011_001101110011 : VALUE=19'b0000000_100011101100;
      15'b011_001101110100 : VALUE=19'b0000000_100011101100;
      15'b011_001101110101 : VALUE=19'b0000000_100011101100;
      15'b011_001101110110 : VALUE=19'b0000000_100011101100;
      15'b011_001101110111 : VALUE=19'b0000000_100011101100;
      15'b011_001101111000 : VALUE=19'b0000000_100011101100;
      15'b011_001101111001 : VALUE=19'b0000000_100011101100;
      15'b011_001101111010 : VALUE=19'b0000000_100011101100;
      15'b011_001101111011 : VALUE=19'b0000000_100011101011;
      15'b011_001101111100 : VALUE=19'b0000000_100011101011;
      15'b011_001101111101 : VALUE=19'b0000000_100011101011;
      15'b011_001101111110 : VALUE=19'b0000000_100011101011;
      15'b011_001101111111 : VALUE=19'b0000000_100011101011;
      15'b011_001110000000 : VALUE=19'b0000000_100011101011;
      15'b011_001110000001 : VALUE=19'b0000000_100011101011;
      15'b011_001110000010 : VALUE=19'b0000000_100011101011;
      15'b011_001110000011 : VALUE=19'b0000000_100011101011;
      15'b011_001110000100 : VALUE=19'b0000000_100011101011;
      15'b011_001110000101 : VALUE=19'b0000000_100011101011;
      15'b011_001110000110 : VALUE=19'b0000000_100011101011;
      15'b011_001110000111 : VALUE=19'b0000000_100011101010;
      15'b011_001110001000 : VALUE=19'b0000000_100011101010;
      15'b011_001110001001 : VALUE=19'b0000000_100011101010;
      15'b011_001110001010 : VALUE=19'b0000000_100011101010;
      15'b011_001110001011 : VALUE=19'b0000000_100011101010;
      15'b011_001110001100 : VALUE=19'b0000000_100011101010;
      15'b011_001110001101 : VALUE=19'b0000000_100011101010;
      15'b011_001110001110 : VALUE=19'b0000000_100011101010;
      15'b011_001110001111 : VALUE=19'b0000000_100011101010;
      15'b011_001110010000 : VALUE=19'b0000000_100011101010;
      15'b011_001110010001 : VALUE=19'b0000000_100011101010;
      15'b011_001110010010 : VALUE=19'b0000000_100011101001;
      15'b011_001110010011 : VALUE=19'b0000000_100011101001;
      15'b011_001110010100 : VALUE=19'b0000000_100011101001;
      15'b011_001110010101 : VALUE=19'b0000000_100011101001;
      15'b011_001110010110 : VALUE=19'b0000000_100011101001;
      15'b011_001110010111 : VALUE=19'b0000000_100011101001;
      15'b011_001110011000 : VALUE=19'b0000000_100011101001;
      15'b011_001110011001 : VALUE=19'b0000000_100011101001;
      15'b011_001110011010 : VALUE=19'b0000000_100011101001;
      15'b011_001110011011 : VALUE=19'b0000000_100011101001;
      15'b011_001110011100 : VALUE=19'b0000000_100011101001;
      15'b011_001110011101 : VALUE=19'b0000000_100011101001;
      15'b011_001110011110 : VALUE=19'b0000000_100011101000;
      15'b011_001110011111 : VALUE=19'b0000000_100011101000;
      15'b011_001110100000 : VALUE=19'b0000000_100011101000;
      15'b011_001110100001 : VALUE=19'b0000000_100011101000;
      15'b011_001110100010 : VALUE=19'b0000000_100011101000;
      15'b011_001110100011 : VALUE=19'b0000000_100011101000;
      15'b011_001110100100 : VALUE=19'b0000000_100011101000;
      15'b011_001110100101 : VALUE=19'b0000000_100011101000;
      15'b011_001110100110 : VALUE=19'b0000000_100011101000;
      15'b011_001110100111 : VALUE=19'b0000000_100011101000;
      15'b011_001110101000 : VALUE=19'b0000000_100011101000;
      15'b011_001110101001 : VALUE=19'b0000000_100011101000;
      15'b011_001110101010 : VALUE=19'b0000000_100011100111;
      15'b011_001110101011 : VALUE=19'b0000000_100011100111;
      15'b011_001110101100 : VALUE=19'b0000000_100011100111;
      15'b011_001110101101 : VALUE=19'b0000000_100011100111;
      15'b011_001110101110 : VALUE=19'b0000000_100011100111;
      15'b011_001110101111 : VALUE=19'b0000000_100011100111;
      15'b011_001110110000 : VALUE=19'b0000000_100011100111;
      15'b011_001110110001 : VALUE=19'b0000000_100011100111;
      15'b011_001110110010 : VALUE=19'b0000000_100011100111;
      15'b011_001110110011 : VALUE=19'b0000000_100011100111;
      15'b011_001110110100 : VALUE=19'b0000000_100011100111;
      15'b011_001110110101 : VALUE=19'b0000000_100011100110;
      15'b011_001110110110 : VALUE=19'b0000000_100011100110;
      15'b011_001110110111 : VALUE=19'b0000000_100011100110;
      15'b011_001110111000 : VALUE=19'b0000000_100011100110;
      15'b011_001110111001 : VALUE=19'b0000000_100011100110;
      15'b011_001110111010 : VALUE=19'b0000000_100011100110;
      15'b011_001110111011 : VALUE=19'b0000000_100011100110;
      15'b011_001110111100 : VALUE=19'b0000000_100011100110;
      15'b011_001110111101 : VALUE=19'b0000000_100011100110;
      15'b011_001110111110 : VALUE=19'b0000000_100011100110;
      15'b011_001110111111 : VALUE=19'b0000000_100011100110;
      15'b011_001111000000 : VALUE=19'b0000000_100011100110;
      15'b011_001111000001 : VALUE=19'b0000000_100011100101;
      15'b011_001111000010 : VALUE=19'b0000000_100011100101;
      15'b011_001111000011 : VALUE=19'b0000000_100011100101;
      15'b011_001111000100 : VALUE=19'b0000000_100011100101;
      15'b011_001111000101 : VALUE=19'b0000000_100011100101;
      15'b011_001111000110 : VALUE=19'b0000000_100011100101;
      15'b011_001111000111 : VALUE=19'b0000000_100011100101;
      15'b011_001111001000 : VALUE=19'b0000000_100011100101;
      15'b011_001111001001 : VALUE=19'b0000000_100011100101;
      15'b011_001111001010 : VALUE=19'b0000000_100011100101;
      15'b011_001111001011 : VALUE=19'b0000000_100011100101;
      15'b011_001111001100 : VALUE=19'b0000000_100011100101;
      15'b011_001111001101 : VALUE=19'b0000000_100011100100;
      15'b011_001111001110 : VALUE=19'b0000000_100011100100;
      15'b011_001111001111 : VALUE=19'b0000000_100011100100;
      15'b011_001111010000 : VALUE=19'b0000000_100011100100;
      15'b011_001111010001 : VALUE=19'b0000000_100011100100;
      15'b011_001111010010 : VALUE=19'b0000000_100011100100;
      15'b011_001111010011 : VALUE=19'b0000000_100011100100;
      15'b011_001111010100 : VALUE=19'b0000000_100011100100;
      15'b011_001111010101 : VALUE=19'b0000000_100011100100;
      15'b011_001111010110 : VALUE=19'b0000000_100011100100;
      15'b011_001111010111 : VALUE=19'b0000000_100011100100;
      15'b011_001111011000 : VALUE=19'b0000000_100011100011;
      15'b011_001111011001 : VALUE=19'b0000000_100011100011;
      15'b011_001111011010 : VALUE=19'b0000000_100011100011;
      15'b011_001111011011 : VALUE=19'b0000000_100011100011;
      15'b011_001111011100 : VALUE=19'b0000000_100011100011;
      15'b011_001111011101 : VALUE=19'b0000000_100011100011;
      15'b011_001111011110 : VALUE=19'b0000000_100011100011;
      15'b011_001111011111 : VALUE=19'b0000000_100011100011;
      15'b011_001111100000 : VALUE=19'b0000000_100011100011;
      15'b011_001111100001 : VALUE=19'b0000000_100011100011;
      15'b011_001111100010 : VALUE=19'b0000000_100011100011;
      15'b011_001111100011 : VALUE=19'b0000000_100011100011;
      15'b011_001111100100 : VALUE=19'b0000000_100011100010;
      15'b011_001111100101 : VALUE=19'b0000000_100011100010;
      15'b011_001111100110 : VALUE=19'b0000000_100011100010;
      15'b011_001111100111 : VALUE=19'b0000000_100011100010;
      15'b011_001111101000 : VALUE=19'b0000000_100011100010;
      15'b011_001111101001 : VALUE=19'b0000000_100011100010;
      15'b011_001111101010 : VALUE=19'b0000000_100011100010;
      15'b011_001111101011 : VALUE=19'b0000000_100011100010;
      15'b011_001111101100 : VALUE=19'b0000000_100011100010;
      15'b011_001111101101 : VALUE=19'b0000000_100011100010;
      15'b011_001111101110 : VALUE=19'b0000000_100011100010;
      15'b011_001111101111 : VALUE=19'b0000000_100011100010;
      15'b011_001111110000 : VALUE=19'b0000000_100011100001;
      15'b011_001111110001 : VALUE=19'b0000000_100011100001;
      15'b011_001111110010 : VALUE=19'b0000000_100011100001;
      15'b011_001111110011 : VALUE=19'b0000000_100011100001;
      15'b011_001111110100 : VALUE=19'b0000000_100011100001;
      15'b011_001111110101 : VALUE=19'b0000000_100011100001;
      15'b011_001111110110 : VALUE=19'b0000000_100011100001;
      15'b011_001111110111 : VALUE=19'b0000000_100011100001;
      15'b011_001111111000 : VALUE=19'b0000000_100011100001;
      15'b011_001111111001 : VALUE=19'b0000000_100011100001;
      15'b011_001111111010 : VALUE=19'b0000000_100011100001;
      15'b011_001111111011 : VALUE=19'b0000000_100011100000;
      15'b011_001111111100 : VALUE=19'b0000000_100011100000;
      15'b011_001111111101 : VALUE=19'b0000000_100011100000;
      15'b011_001111111110 : VALUE=19'b0000000_100011100000;
      15'b011_001111111111 : VALUE=19'b0000000_100011100000;
      15'b011_010000000000 : VALUE=19'b0000000_100011100000;
      15'b011_010000000001 : VALUE=19'b0000000_100011100000;
      15'b011_010000000010 : VALUE=19'b0000000_100011100000;
      15'b011_010000000011 : VALUE=19'b0000000_100011100000;
      15'b011_010000000100 : VALUE=19'b0000000_100011100000;
      15'b011_010000000101 : VALUE=19'b0000000_100011100000;
      15'b011_010000000110 : VALUE=19'b0000000_100011100000;
      15'b011_010000000111 : VALUE=19'b0000000_100011011111;
      15'b011_010000001000 : VALUE=19'b0000000_100011011111;
      15'b011_010000001001 : VALUE=19'b0000000_100011011111;
      15'b011_010000001010 : VALUE=19'b0000000_100011011111;
      15'b011_010000001011 : VALUE=19'b0000000_100011011111;
      15'b011_010000001100 : VALUE=19'b0000000_100011011111;
      15'b011_010000001101 : VALUE=19'b0000000_100011011111;
      15'b011_010000001110 : VALUE=19'b0000000_100011011111;
      15'b011_010000001111 : VALUE=19'b0000000_100011011111;
      15'b011_010000010000 : VALUE=19'b0000000_100011011111;
      15'b011_010000010001 : VALUE=19'b0000000_100011011111;
      15'b011_010000010010 : VALUE=19'b0000000_100011011111;
      15'b011_010000010011 : VALUE=19'b0000000_100011011110;
      15'b011_010000010100 : VALUE=19'b0000000_100011011110;
      15'b011_010000010101 : VALUE=19'b0000000_100011011110;
      15'b011_010000010110 : VALUE=19'b0000000_100011011110;
      15'b011_010000010111 : VALUE=19'b0000000_100011011110;
      15'b011_010000011000 : VALUE=19'b0000000_100011011110;
      15'b011_010000011001 : VALUE=19'b0000000_100011011110;
      15'b011_010000011010 : VALUE=19'b0000000_100011011110;
      15'b011_010000011011 : VALUE=19'b0000000_100011011110;
      15'b011_010000011100 : VALUE=19'b0000000_100011011110;
      15'b011_010000011101 : VALUE=19'b0000000_100011011110;
      15'b011_010000011110 : VALUE=19'b0000000_100011011101;
      15'b011_010000011111 : VALUE=19'b0000000_100011011101;
      15'b011_010000100000 : VALUE=19'b0000000_100011011101;
      15'b011_010000100001 : VALUE=19'b0000000_100011011101;
      15'b011_010000100010 : VALUE=19'b0000000_100011011101;
      15'b011_010000100011 : VALUE=19'b0000000_100011011101;
      15'b011_010000100100 : VALUE=19'b0000000_100011011101;
      15'b011_010000100101 : VALUE=19'b0000000_100011011101;
      15'b011_010000100110 : VALUE=19'b0000000_100011011101;
      15'b011_010000100111 : VALUE=19'b0000000_100011011101;
      15'b011_010000101000 : VALUE=19'b0000000_100011011101;
      15'b011_010000101001 : VALUE=19'b0000000_100011011101;
      15'b011_010000101010 : VALUE=19'b0000000_100011011100;
      15'b011_010000101011 : VALUE=19'b0000000_100011011100;
      15'b011_010000101100 : VALUE=19'b0000000_100011011100;
      15'b011_010000101101 : VALUE=19'b0000000_100011011100;
      15'b011_010000101110 : VALUE=19'b0000000_100011011100;
      15'b011_010000101111 : VALUE=19'b0000000_100011011100;
      15'b011_010000110000 : VALUE=19'b0000000_100011011100;
      15'b011_010000110001 : VALUE=19'b0000000_100011011100;
      15'b011_010000110010 : VALUE=19'b0000000_100011011100;
      15'b011_010000110011 : VALUE=19'b0000000_100011011100;
      15'b011_010000110100 : VALUE=19'b0000000_100011011100;
      15'b011_010000110101 : VALUE=19'b0000000_100011011100;
      15'b011_010000110110 : VALUE=19'b0000000_100011011011;
      15'b011_010000110111 : VALUE=19'b0000000_100011011011;
      15'b011_010000111000 : VALUE=19'b0000000_100011011011;
      15'b011_010000111001 : VALUE=19'b0000000_100011011011;
      15'b011_010000111010 : VALUE=19'b0000000_100011011011;
      15'b011_010000111011 : VALUE=19'b0000000_100011011011;
      15'b011_010000111100 : VALUE=19'b0000000_100011011011;
      15'b011_010000111101 : VALUE=19'b0000000_100011011011;
      15'b011_010000111110 : VALUE=19'b0000000_100011011011;
      15'b011_010000111111 : VALUE=19'b0000000_100011011011;
      15'b011_010001000000 : VALUE=19'b0000000_100011011011;
      15'b011_010001000001 : VALUE=19'b0000000_100011011011;
      15'b011_010001000010 : VALUE=19'b0000000_100011011010;
      15'b011_010001000011 : VALUE=19'b0000000_100011011010;
      15'b011_010001000100 : VALUE=19'b0000000_100011011010;
      15'b011_010001000101 : VALUE=19'b0000000_100011011010;
      15'b011_010001000110 : VALUE=19'b0000000_100011011010;
      15'b011_010001000111 : VALUE=19'b0000000_100011011010;
      15'b011_010001001000 : VALUE=19'b0000000_100011011010;
      15'b011_010001001001 : VALUE=19'b0000000_100011011010;
      15'b011_010001001010 : VALUE=19'b0000000_100011011010;
      15'b011_010001001011 : VALUE=19'b0000000_100011011010;
      15'b011_010001001100 : VALUE=19'b0000000_100011011010;
      15'b011_010001001101 : VALUE=19'b0000000_100011011010;
      15'b011_010001001110 : VALUE=19'b0000000_100011011001;
      15'b011_010001001111 : VALUE=19'b0000000_100011011001;
      15'b011_010001010000 : VALUE=19'b0000000_100011011001;
      15'b011_010001010001 : VALUE=19'b0000000_100011011001;
      15'b011_010001010010 : VALUE=19'b0000000_100011011001;
      15'b011_010001010011 : VALUE=19'b0000000_100011011001;
      15'b011_010001010100 : VALUE=19'b0000000_100011011001;
      15'b011_010001010101 : VALUE=19'b0000000_100011011001;
      15'b011_010001010110 : VALUE=19'b0000000_100011011001;
      15'b011_010001010111 : VALUE=19'b0000000_100011011001;
      15'b011_010001011000 : VALUE=19'b0000000_100011011001;
      15'b011_010001011001 : VALUE=19'b0000000_100011011000;
      15'b011_010001011010 : VALUE=19'b0000000_100011011000;
      15'b011_010001011011 : VALUE=19'b0000000_100011011000;
      15'b011_010001011100 : VALUE=19'b0000000_100011011000;
      15'b011_010001011101 : VALUE=19'b0000000_100011011000;
      15'b011_010001011110 : VALUE=19'b0000000_100011011000;
      15'b011_010001011111 : VALUE=19'b0000000_100011011000;
      15'b011_010001100000 : VALUE=19'b0000000_100011011000;
      15'b011_010001100001 : VALUE=19'b0000000_100011011000;
      15'b011_010001100010 : VALUE=19'b0000000_100011011000;
      15'b011_010001100011 : VALUE=19'b0000000_100011011000;
      15'b011_010001100100 : VALUE=19'b0000000_100011011000;
      15'b011_010001100101 : VALUE=19'b0000000_100011010111;
      15'b011_010001100110 : VALUE=19'b0000000_100011010111;
      15'b011_010001100111 : VALUE=19'b0000000_100011010111;
      15'b011_010001101000 : VALUE=19'b0000000_100011010111;
      15'b011_010001101001 : VALUE=19'b0000000_100011010111;
      15'b011_010001101010 : VALUE=19'b0000000_100011010111;
      15'b011_010001101011 : VALUE=19'b0000000_100011010111;
      15'b011_010001101100 : VALUE=19'b0000000_100011010111;
      15'b011_010001101101 : VALUE=19'b0000000_100011010111;
      15'b011_010001101110 : VALUE=19'b0000000_100011010111;
      15'b011_010001101111 : VALUE=19'b0000000_100011010111;
      15'b011_010001110000 : VALUE=19'b0000000_100011010111;
      15'b011_010001110001 : VALUE=19'b0000000_100011010110;
      15'b011_010001110010 : VALUE=19'b0000000_100011010110;
      15'b011_010001110011 : VALUE=19'b0000000_100011010110;
      15'b011_010001110100 : VALUE=19'b0000000_100011010110;
      15'b011_010001110101 : VALUE=19'b0000000_100011010110;
      15'b011_010001110110 : VALUE=19'b0000000_100011010110;
      15'b011_010001110111 : VALUE=19'b0000000_100011010110;
      15'b011_010001111000 : VALUE=19'b0000000_100011010110;
      15'b011_010001111001 : VALUE=19'b0000000_100011010110;
      15'b011_010001111010 : VALUE=19'b0000000_100011010110;
      15'b011_010001111011 : VALUE=19'b0000000_100011010110;
      15'b011_010001111100 : VALUE=19'b0000000_100011010110;
      15'b011_010001111101 : VALUE=19'b0000000_100011010101;
      15'b011_010001111110 : VALUE=19'b0000000_100011010101;
      15'b011_010001111111 : VALUE=19'b0000000_100011010101;
      15'b011_010010000000 : VALUE=19'b0000000_100011010101;
      15'b011_010010000001 : VALUE=19'b0000000_100011010101;
      15'b011_010010000010 : VALUE=19'b0000000_100011010101;
      15'b011_010010000011 : VALUE=19'b0000000_100011010101;
      15'b011_010010000100 : VALUE=19'b0000000_100011010101;
      15'b011_010010000101 : VALUE=19'b0000000_100011010101;
      15'b011_010010000110 : VALUE=19'b0000000_100011010101;
      15'b011_010010000111 : VALUE=19'b0000000_100011010101;
      15'b011_010010001000 : VALUE=19'b0000000_100011010101;
      15'b011_010010001001 : VALUE=19'b0000000_100011010100;
      15'b011_010010001010 : VALUE=19'b0000000_100011010100;
      15'b011_010010001011 : VALUE=19'b0000000_100011010100;
      15'b011_010010001100 : VALUE=19'b0000000_100011010100;
      15'b011_010010001101 : VALUE=19'b0000000_100011010100;
      15'b011_010010001110 : VALUE=19'b0000000_100011010100;
      15'b011_010010001111 : VALUE=19'b0000000_100011010100;
      15'b011_010010010000 : VALUE=19'b0000000_100011010100;
      15'b011_010010010001 : VALUE=19'b0000000_100011010100;
      15'b011_010010010010 : VALUE=19'b0000000_100011010100;
      15'b011_010010010011 : VALUE=19'b0000000_100011010100;
      15'b011_010010010100 : VALUE=19'b0000000_100011010100;
      15'b011_010010010101 : VALUE=19'b0000000_100011010011;
      15'b011_010010010110 : VALUE=19'b0000000_100011010011;
      15'b011_010010010111 : VALUE=19'b0000000_100011010011;
      15'b011_010010011000 : VALUE=19'b0000000_100011010011;
      15'b011_010010011001 : VALUE=19'b0000000_100011010011;
      15'b011_010010011010 : VALUE=19'b0000000_100011010011;
      15'b011_010010011011 : VALUE=19'b0000000_100011010011;
      15'b011_010010011100 : VALUE=19'b0000000_100011010011;
      15'b011_010010011101 : VALUE=19'b0000000_100011010011;
      15'b011_010010011110 : VALUE=19'b0000000_100011010011;
      15'b011_010010011111 : VALUE=19'b0000000_100011010011;
      15'b011_010010100000 : VALUE=19'b0000000_100011010011;
      15'b011_010010100001 : VALUE=19'b0000000_100011010010;
      15'b011_010010100010 : VALUE=19'b0000000_100011010010;
      15'b011_010010100011 : VALUE=19'b0000000_100011010010;
      15'b011_010010100100 : VALUE=19'b0000000_100011010010;
      15'b011_010010100101 : VALUE=19'b0000000_100011010010;
      15'b011_010010100110 : VALUE=19'b0000000_100011010010;
      15'b011_010010100111 : VALUE=19'b0000000_100011010010;
      15'b011_010010101000 : VALUE=19'b0000000_100011010010;
      15'b011_010010101001 : VALUE=19'b0000000_100011010010;
      15'b011_010010101010 : VALUE=19'b0000000_100011010010;
      15'b011_010010101011 : VALUE=19'b0000000_100011010010;
      15'b011_010010101100 : VALUE=19'b0000000_100011010010;
      15'b011_010010101101 : VALUE=19'b0000000_100011010001;
      15'b011_010010101110 : VALUE=19'b0000000_100011010001;
      15'b011_010010101111 : VALUE=19'b0000000_100011010001;
      15'b011_010010110000 : VALUE=19'b0000000_100011010001;
      15'b011_010010110001 : VALUE=19'b0000000_100011010001;
      15'b011_010010110010 : VALUE=19'b0000000_100011010001;
      15'b011_010010110011 : VALUE=19'b0000000_100011010001;
      15'b011_010010110100 : VALUE=19'b0000000_100011010001;
      15'b011_010010110101 : VALUE=19'b0000000_100011010001;
      15'b011_010010110110 : VALUE=19'b0000000_100011010001;
      15'b011_010010110111 : VALUE=19'b0000000_100011010001;
      15'b011_010010111000 : VALUE=19'b0000000_100011010001;
      15'b011_010010111001 : VALUE=19'b0000000_100011010000;
      15'b011_010010111010 : VALUE=19'b0000000_100011010000;
      15'b011_010010111011 : VALUE=19'b0000000_100011010000;
      15'b011_010010111100 : VALUE=19'b0000000_100011010000;
      15'b011_010010111101 : VALUE=19'b0000000_100011010000;
      15'b011_010010111110 : VALUE=19'b0000000_100011010000;
      15'b011_010010111111 : VALUE=19'b0000000_100011010000;
      15'b011_010011000000 : VALUE=19'b0000000_100011010000;
      15'b011_010011000001 : VALUE=19'b0000000_100011010000;
      15'b011_010011000010 : VALUE=19'b0000000_100011010000;
      15'b011_010011000011 : VALUE=19'b0000000_100011010000;
      15'b011_010011000100 : VALUE=19'b0000000_100011010000;
      15'b011_010011000101 : VALUE=19'b0000000_100011001111;
      15'b011_010011000110 : VALUE=19'b0000000_100011001111;
      15'b011_010011000111 : VALUE=19'b0000000_100011001111;
      15'b011_010011001000 : VALUE=19'b0000000_100011001111;
      15'b011_010011001001 : VALUE=19'b0000000_100011001111;
      15'b011_010011001010 : VALUE=19'b0000000_100011001111;
      15'b011_010011001011 : VALUE=19'b0000000_100011001111;
      15'b011_010011001100 : VALUE=19'b0000000_100011001111;
      15'b011_010011001101 : VALUE=19'b0000000_100011001111;
      15'b011_010011001110 : VALUE=19'b0000000_100011001111;
      15'b011_010011001111 : VALUE=19'b0000000_100011001111;
      15'b011_010011010000 : VALUE=19'b0000000_100011001111;
      15'b011_010011010001 : VALUE=19'b0000000_100011001110;
      15'b011_010011010010 : VALUE=19'b0000000_100011001110;
      15'b011_010011010011 : VALUE=19'b0000000_100011001110;
      15'b011_010011010100 : VALUE=19'b0000000_100011001110;
      15'b011_010011010101 : VALUE=19'b0000000_100011001110;
      15'b011_010011010110 : VALUE=19'b0000000_100011001110;
      15'b011_010011010111 : VALUE=19'b0000000_100011001110;
      15'b011_010011011000 : VALUE=19'b0000000_100011001110;
      15'b011_010011011001 : VALUE=19'b0000000_100011001110;
      15'b011_010011011010 : VALUE=19'b0000000_100011001110;
      15'b011_010011011011 : VALUE=19'b0000000_100011001110;
      15'b011_010011011100 : VALUE=19'b0000000_100011001110;
      15'b011_010011011101 : VALUE=19'b0000000_100011001101;
      15'b011_010011011110 : VALUE=19'b0000000_100011001101;
      15'b011_010011011111 : VALUE=19'b0000000_100011001101;
      15'b011_010011100000 : VALUE=19'b0000000_100011001101;
      15'b011_010011100001 : VALUE=19'b0000000_100011001101;
      15'b011_010011100010 : VALUE=19'b0000000_100011001101;
      15'b011_010011100011 : VALUE=19'b0000000_100011001101;
      15'b011_010011100100 : VALUE=19'b0000000_100011001101;
      15'b011_010011100101 : VALUE=19'b0000000_100011001101;
      15'b011_010011100110 : VALUE=19'b0000000_100011001101;
      15'b011_010011100111 : VALUE=19'b0000000_100011001101;
      15'b011_010011101000 : VALUE=19'b0000000_100011001101;
      15'b011_010011101001 : VALUE=19'b0000000_100011001100;
      15'b011_010011101010 : VALUE=19'b0000000_100011001100;
      15'b011_010011101011 : VALUE=19'b0000000_100011001100;
      15'b011_010011101100 : VALUE=19'b0000000_100011001100;
      15'b011_010011101101 : VALUE=19'b0000000_100011001100;
      15'b011_010011101110 : VALUE=19'b0000000_100011001100;
      15'b011_010011101111 : VALUE=19'b0000000_100011001100;
      15'b011_010011110000 : VALUE=19'b0000000_100011001100;
      15'b011_010011110001 : VALUE=19'b0000000_100011001100;
      15'b011_010011110010 : VALUE=19'b0000000_100011001100;
      15'b011_010011110011 : VALUE=19'b0000000_100011001100;
      15'b011_010011110100 : VALUE=19'b0000000_100011001100;
      15'b011_010011110101 : VALUE=19'b0000000_100011001011;
      15'b011_010011110110 : VALUE=19'b0000000_100011001011;
      15'b011_010011110111 : VALUE=19'b0000000_100011001011;
      15'b011_010011111000 : VALUE=19'b0000000_100011001011;
      15'b011_010011111001 : VALUE=19'b0000000_100011001011;
      15'b011_010011111010 : VALUE=19'b0000000_100011001011;
      15'b011_010011111011 : VALUE=19'b0000000_100011001011;
      15'b011_010011111100 : VALUE=19'b0000000_100011001011;
      15'b011_010011111101 : VALUE=19'b0000000_100011001011;
      15'b011_010011111110 : VALUE=19'b0000000_100011001011;
      15'b011_010011111111 : VALUE=19'b0000000_100011001011;
      15'b011_010100000000 : VALUE=19'b0000000_100011001011;
      15'b011_010100000001 : VALUE=19'b0000000_100011001010;
      15'b011_010100000010 : VALUE=19'b0000000_100011001010;
      15'b011_010100000011 : VALUE=19'b0000000_100011001010;
      15'b011_010100000100 : VALUE=19'b0000000_100011001010;
      15'b011_010100000101 : VALUE=19'b0000000_100011001010;
      15'b011_010100000110 : VALUE=19'b0000000_100011001010;
      15'b011_010100000111 : VALUE=19'b0000000_100011001010;
      15'b011_010100001000 : VALUE=19'b0000000_100011001010;
      15'b011_010100001001 : VALUE=19'b0000000_100011001010;
      15'b011_010100001010 : VALUE=19'b0000000_100011001010;
      15'b011_010100001011 : VALUE=19'b0000000_100011001010;
      15'b011_010100001100 : VALUE=19'b0000000_100011001010;
      15'b011_010100001101 : VALUE=19'b0000000_100011001001;
      15'b011_010100001110 : VALUE=19'b0000000_100011001001;
      15'b011_010100001111 : VALUE=19'b0000000_100011001001;
      15'b011_010100010000 : VALUE=19'b0000000_100011001001;
      15'b011_010100010001 : VALUE=19'b0000000_100011001001;
      15'b011_010100010010 : VALUE=19'b0000000_100011001001;
      15'b011_010100010011 : VALUE=19'b0000000_100011001001;
      15'b011_010100010100 : VALUE=19'b0000000_100011001001;
      15'b011_010100010101 : VALUE=19'b0000000_100011001001;
      15'b011_010100010110 : VALUE=19'b0000000_100011001001;
      15'b011_010100010111 : VALUE=19'b0000000_100011001001;
      15'b011_010100011000 : VALUE=19'b0000000_100011001001;
      15'b011_010100011001 : VALUE=19'b0000000_100011001000;
      15'b011_010100011010 : VALUE=19'b0000000_100011001000;
      15'b011_010100011011 : VALUE=19'b0000000_100011001000;
      15'b011_010100011100 : VALUE=19'b0000000_100011001000;
      15'b011_010100011101 : VALUE=19'b0000000_100011001000;
      15'b011_010100011110 : VALUE=19'b0000000_100011001000;
      15'b011_010100011111 : VALUE=19'b0000000_100011001000;
      15'b011_010100100000 : VALUE=19'b0000000_100011001000;
      15'b011_010100100001 : VALUE=19'b0000000_100011001000;
      15'b011_010100100010 : VALUE=19'b0000000_100011001000;
      15'b011_010100100011 : VALUE=19'b0000000_100011001000;
      15'b011_010100100100 : VALUE=19'b0000000_100011001000;
      15'b011_010100100101 : VALUE=19'b0000000_100011000111;
      15'b011_010100100110 : VALUE=19'b0000000_100011000111;
      15'b011_010100100111 : VALUE=19'b0000000_100011000111;
      15'b011_010100101000 : VALUE=19'b0000000_100011000111;
      15'b011_010100101001 : VALUE=19'b0000000_100011000111;
      15'b011_010100101010 : VALUE=19'b0000000_100011000111;
      15'b011_010100101011 : VALUE=19'b0000000_100011000111;
      15'b011_010100101100 : VALUE=19'b0000000_100011000111;
      15'b011_010100101101 : VALUE=19'b0000000_100011000111;
      15'b011_010100101110 : VALUE=19'b0000000_100011000111;
      15'b011_010100101111 : VALUE=19'b0000000_100011000111;
      15'b011_010100110000 : VALUE=19'b0000000_100011000111;
      15'b011_010100110001 : VALUE=19'b0000000_100011000110;
      15'b011_010100110010 : VALUE=19'b0000000_100011000110;
      15'b011_010100110011 : VALUE=19'b0000000_100011000110;
      15'b011_010100110100 : VALUE=19'b0000000_100011000110;
      15'b011_010100110101 : VALUE=19'b0000000_100011000110;
      15'b011_010100110110 : VALUE=19'b0000000_100011000110;
      15'b011_010100110111 : VALUE=19'b0000000_100011000110;
      15'b011_010100111000 : VALUE=19'b0000000_100011000110;
      15'b011_010100111001 : VALUE=19'b0000000_100011000110;
      15'b011_010100111010 : VALUE=19'b0000000_100011000110;
      15'b011_010100111011 : VALUE=19'b0000000_100011000110;
      15'b011_010100111100 : VALUE=19'b0000000_100011000110;
      15'b011_010100111101 : VALUE=19'b0000000_100011000101;
      15'b011_010100111110 : VALUE=19'b0000000_100011000101;
      15'b011_010100111111 : VALUE=19'b0000000_100011000101;
      15'b011_010101000000 : VALUE=19'b0000000_100011000101;
      15'b011_010101000001 : VALUE=19'b0000000_100011000101;
      15'b011_010101000010 : VALUE=19'b0000000_100011000101;
      15'b011_010101000011 : VALUE=19'b0000000_100011000101;
      15'b011_010101000100 : VALUE=19'b0000000_100011000101;
      15'b011_010101000101 : VALUE=19'b0000000_100011000101;
      15'b011_010101000110 : VALUE=19'b0000000_100011000101;
      15'b011_010101000111 : VALUE=19'b0000000_100011000101;
      15'b011_010101001000 : VALUE=19'b0000000_100011000101;
      15'b011_010101001001 : VALUE=19'b0000000_100011000100;
      15'b011_010101001010 : VALUE=19'b0000000_100011000100;
      15'b011_010101001011 : VALUE=19'b0000000_100011000100;
      15'b011_010101001100 : VALUE=19'b0000000_100011000100;
      15'b011_010101001101 : VALUE=19'b0000000_100011000100;
      15'b011_010101001110 : VALUE=19'b0000000_100011000100;
      15'b011_010101001111 : VALUE=19'b0000000_100011000100;
      15'b011_010101010000 : VALUE=19'b0000000_100011000100;
      15'b011_010101010001 : VALUE=19'b0000000_100011000100;
      15'b011_010101010010 : VALUE=19'b0000000_100011000100;
      15'b011_010101010011 : VALUE=19'b0000000_100011000100;
      15'b011_010101010100 : VALUE=19'b0000000_100011000100;
      15'b011_010101010101 : VALUE=19'b0000000_100011000011;
      15'b011_010101010110 : VALUE=19'b0000000_100011000011;
      15'b011_010101010111 : VALUE=19'b0000000_100011000011;
      15'b011_010101011000 : VALUE=19'b0000000_100011000011;
      15'b011_010101011001 : VALUE=19'b0000000_100011000011;
      15'b011_010101011010 : VALUE=19'b0000000_100011000011;
      15'b011_010101011011 : VALUE=19'b0000000_100011000011;
      15'b011_010101011100 : VALUE=19'b0000000_100011000011;
      15'b011_010101011101 : VALUE=19'b0000000_100011000011;
      15'b011_010101011110 : VALUE=19'b0000000_100011000011;
      15'b011_010101011111 : VALUE=19'b0000000_100011000011;
      15'b011_010101100000 : VALUE=19'b0000000_100011000011;
      15'b011_010101100001 : VALUE=19'b0000000_100011000011;
      15'b011_010101100010 : VALUE=19'b0000000_100011000010;
      15'b011_010101100011 : VALUE=19'b0000000_100011000010;
      15'b011_010101100100 : VALUE=19'b0000000_100011000010;
      15'b011_010101100101 : VALUE=19'b0000000_100011000010;
      15'b011_010101100110 : VALUE=19'b0000000_100011000010;
      15'b011_010101100111 : VALUE=19'b0000000_100011000010;
      15'b011_010101101000 : VALUE=19'b0000000_100011000010;
      15'b011_010101101001 : VALUE=19'b0000000_100011000010;
      15'b011_010101101010 : VALUE=19'b0000000_100011000010;
      15'b011_010101101011 : VALUE=19'b0000000_100011000010;
      15'b011_010101101100 : VALUE=19'b0000000_100011000010;
      15'b011_010101101101 : VALUE=19'b0000000_100011000010;
      15'b011_010101101110 : VALUE=19'b0000000_100011000001;
      15'b011_010101101111 : VALUE=19'b0000000_100011000001;
      15'b011_010101110000 : VALUE=19'b0000000_100011000001;
      15'b011_010101110001 : VALUE=19'b0000000_100011000001;
      15'b011_010101110010 : VALUE=19'b0000000_100011000001;
      15'b011_010101110011 : VALUE=19'b0000000_100011000001;
      15'b011_010101110100 : VALUE=19'b0000000_100011000001;
      15'b011_010101110101 : VALUE=19'b0000000_100011000001;
      15'b011_010101110110 : VALUE=19'b0000000_100011000001;
      15'b011_010101110111 : VALUE=19'b0000000_100011000001;
      15'b011_010101111000 : VALUE=19'b0000000_100011000001;
      15'b011_010101111001 : VALUE=19'b0000000_100011000001;
      15'b011_010101111010 : VALUE=19'b0000000_100011000000;
      15'b011_010101111011 : VALUE=19'b0000000_100011000000;
      15'b011_010101111100 : VALUE=19'b0000000_100011000000;
      15'b011_010101111101 : VALUE=19'b0000000_100011000000;
      15'b011_010101111110 : VALUE=19'b0000000_100011000000;
      15'b011_010101111111 : VALUE=19'b0000000_100011000000;
      15'b011_010110000000 : VALUE=19'b0000000_100011000000;
      15'b011_010110000001 : VALUE=19'b0000000_100011000000;
      15'b011_010110000010 : VALUE=19'b0000000_100011000000;
      15'b011_010110000011 : VALUE=19'b0000000_100011000000;
      15'b011_010110000100 : VALUE=19'b0000000_100011000000;
      15'b011_010110000101 : VALUE=19'b0000000_100011000000;
      15'b011_010110000110 : VALUE=19'b0000000_100010111111;
      15'b011_010110000111 : VALUE=19'b0000000_100010111111;
      15'b011_010110001000 : VALUE=19'b0000000_100010111111;
      15'b011_010110001001 : VALUE=19'b0000000_100010111111;
      15'b011_010110001010 : VALUE=19'b0000000_100010111111;
      15'b011_010110001011 : VALUE=19'b0000000_100010111111;
      15'b011_010110001100 : VALUE=19'b0000000_100010111111;
      15'b011_010110001101 : VALUE=19'b0000000_100010111111;
      15'b011_010110001110 : VALUE=19'b0000000_100010111111;
      15'b011_010110001111 : VALUE=19'b0000000_100010111111;
      15'b011_010110010000 : VALUE=19'b0000000_100010111111;
      15'b011_010110010001 : VALUE=19'b0000000_100010111111;
      15'b011_010110010010 : VALUE=19'b0000000_100010111111;
      15'b011_010110010011 : VALUE=19'b0000000_100010111110;
      15'b011_010110010100 : VALUE=19'b0000000_100010111110;
      15'b011_010110010101 : VALUE=19'b0000000_100010111110;
      15'b011_010110010110 : VALUE=19'b0000000_100010111110;
      15'b011_010110010111 : VALUE=19'b0000000_100010111110;
      15'b011_010110011000 : VALUE=19'b0000000_100010111110;
      15'b011_010110011001 : VALUE=19'b0000000_100010111110;
      15'b011_010110011010 : VALUE=19'b0000000_100010111110;
      15'b011_010110011011 : VALUE=19'b0000000_100010111110;
      15'b011_010110011100 : VALUE=19'b0000000_100010111110;
      15'b011_010110011101 : VALUE=19'b0000000_100010111110;
      15'b011_010110011110 : VALUE=19'b0000000_100010111110;
      15'b011_010110011111 : VALUE=19'b0000000_100010111101;
      15'b011_010110100000 : VALUE=19'b0000000_100010111101;
      15'b011_010110100001 : VALUE=19'b0000000_100010111101;
      15'b011_010110100010 : VALUE=19'b0000000_100010111101;
      15'b011_010110100011 : VALUE=19'b0000000_100010111101;
      15'b011_010110100100 : VALUE=19'b0000000_100010111101;
      15'b011_010110100101 : VALUE=19'b0000000_100010111101;
      15'b011_010110100110 : VALUE=19'b0000000_100010111101;
      15'b011_010110100111 : VALUE=19'b0000000_100010111101;
      15'b011_010110101000 : VALUE=19'b0000000_100010111101;
      15'b011_010110101001 : VALUE=19'b0000000_100010111101;
      15'b011_010110101010 : VALUE=19'b0000000_100010111101;
      15'b011_010110101011 : VALUE=19'b0000000_100010111100;
      15'b011_010110101100 : VALUE=19'b0000000_100010111100;
      15'b011_010110101101 : VALUE=19'b0000000_100010111100;
      15'b011_010110101110 : VALUE=19'b0000000_100010111100;
      15'b011_010110101111 : VALUE=19'b0000000_100010111100;
      15'b011_010110110000 : VALUE=19'b0000000_100010111100;
      15'b011_010110110001 : VALUE=19'b0000000_100010111100;
      15'b011_010110110010 : VALUE=19'b0000000_100010111100;
      15'b011_010110110011 : VALUE=19'b0000000_100010111100;
      15'b011_010110110100 : VALUE=19'b0000000_100010111100;
      15'b011_010110110101 : VALUE=19'b0000000_100010111100;
      15'b011_010110110110 : VALUE=19'b0000000_100010111100;
      15'b011_010110110111 : VALUE=19'b0000000_100010111011;
      15'b011_010110111000 : VALUE=19'b0000000_100010111011;
      15'b011_010110111001 : VALUE=19'b0000000_100010111011;
      15'b011_010110111010 : VALUE=19'b0000000_100010111011;
      15'b011_010110111011 : VALUE=19'b0000000_100010111011;
      15'b011_010110111100 : VALUE=19'b0000000_100010111011;
      15'b011_010110111101 : VALUE=19'b0000000_100010111011;
      15'b011_010110111110 : VALUE=19'b0000000_100010111011;
      15'b011_010110111111 : VALUE=19'b0000000_100010111011;
      15'b011_010111000000 : VALUE=19'b0000000_100010111011;
      15'b011_010111000001 : VALUE=19'b0000000_100010111011;
      15'b011_010111000010 : VALUE=19'b0000000_100010111011;
      15'b011_010111000011 : VALUE=19'b0000000_100010111011;
      15'b011_010111000100 : VALUE=19'b0000000_100010111010;
      15'b011_010111000101 : VALUE=19'b0000000_100010111010;
      15'b011_010111000110 : VALUE=19'b0000000_100010111010;
      15'b011_010111000111 : VALUE=19'b0000000_100010111010;
      15'b011_010111001000 : VALUE=19'b0000000_100010111010;
      15'b011_010111001001 : VALUE=19'b0000000_100010111010;
      15'b011_010111001010 : VALUE=19'b0000000_100010111010;
      15'b011_010111001011 : VALUE=19'b0000000_100010111010;
      15'b011_010111001100 : VALUE=19'b0000000_100010111010;
      15'b011_010111001101 : VALUE=19'b0000000_100010111010;
      15'b011_010111001110 : VALUE=19'b0000000_100010111010;
      15'b011_010111001111 : VALUE=19'b0000000_100010111010;
      15'b011_010111010000 : VALUE=19'b0000000_100010111001;
      15'b011_010111010001 : VALUE=19'b0000000_100010111001;
      15'b011_010111010010 : VALUE=19'b0000000_100010111001;
      15'b011_010111010011 : VALUE=19'b0000000_100010111001;
      15'b011_010111010100 : VALUE=19'b0000000_100010111001;
      15'b011_010111010101 : VALUE=19'b0000000_100010111001;
      15'b011_010111010110 : VALUE=19'b0000000_100010111001;
      15'b011_010111010111 : VALUE=19'b0000000_100010111001;
      15'b011_010111011000 : VALUE=19'b0000000_100010111001;
      15'b011_010111011001 : VALUE=19'b0000000_100010111001;
      15'b011_010111011010 : VALUE=19'b0000000_100010111001;
      15'b011_010111011011 : VALUE=19'b0000000_100010111001;
      15'b011_010111011100 : VALUE=19'b0000000_100010111000;
      15'b011_010111011101 : VALUE=19'b0000000_100010111000;
      15'b011_010111011110 : VALUE=19'b0000000_100010111000;
      15'b011_010111011111 : VALUE=19'b0000000_100010111000;
      15'b011_010111100000 : VALUE=19'b0000000_100010111000;
      15'b011_010111100001 : VALUE=19'b0000000_100010111000;
      15'b011_010111100010 : VALUE=19'b0000000_100010111000;
      15'b011_010111100011 : VALUE=19'b0000000_100010111000;
      15'b011_010111100100 : VALUE=19'b0000000_100010111000;
      15'b011_010111100101 : VALUE=19'b0000000_100010111000;
      15'b011_010111100110 : VALUE=19'b0000000_100010111000;
      15'b011_010111100111 : VALUE=19'b0000000_100010111000;
      15'b011_010111101000 : VALUE=19'b0000000_100010111000;
      15'b011_010111101001 : VALUE=19'b0000000_100010110111;
      15'b011_010111101010 : VALUE=19'b0000000_100010110111;
      15'b011_010111101011 : VALUE=19'b0000000_100010110111;
      15'b011_010111101100 : VALUE=19'b0000000_100010110111;
      15'b011_010111101101 : VALUE=19'b0000000_100010110111;
      15'b011_010111101110 : VALUE=19'b0000000_100010110111;
      15'b011_010111101111 : VALUE=19'b0000000_100010110111;
      15'b011_010111110000 : VALUE=19'b0000000_100010110111;
      15'b011_010111110001 : VALUE=19'b0000000_100010110111;
      15'b011_010111110010 : VALUE=19'b0000000_100010110111;
      15'b011_010111110011 : VALUE=19'b0000000_100010110111;
      15'b011_010111110100 : VALUE=19'b0000000_100010110111;
      15'b011_010111110101 : VALUE=19'b0000000_100010110110;
      15'b011_010111110110 : VALUE=19'b0000000_100010110110;
      15'b011_010111110111 : VALUE=19'b0000000_100010110110;
      15'b011_010111111000 : VALUE=19'b0000000_100010110110;
      15'b011_010111111001 : VALUE=19'b0000000_100010110110;
      15'b011_010111111010 : VALUE=19'b0000000_100010110110;
      15'b011_010111111011 : VALUE=19'b0000000_100010110110;
      15'b011_010111111100 : VALUE=19'b0000000_100010110110;
      15'b011_010111111101 : VALUE=19'b0000000_100010110110;
      15'b011_010111111110 : VALUE=19'b0000000_100010110110;
      15'b011_010111111111 : VALUE=19'b0000000_100010110110;
      15'b011_011000000000 : VALUE=19'b0000000_100010110110;
      15'b011_011000000001 : VALUE=19'b0000000_100010110101;
      15'b011_011000000010 : VALUE=19'b0000000_100010110101;
      15'b011_011000000011 : VALUE=19'b0000000_100010110101;
      15'b011_011000000100 : VALUE=19'b0000000_100010110101;
      15'b011_011000000101 : VALUE=19'b0000000_100010110101;
      15'b011_011000000110 : VALUE=19'b0000000_100010110101;
      15'b011_011000000111 : VALUE=19'b0000000_100010110101;
      15'b011_011000001000 : VALUE=19'b0000000_100010110101;
      15'b011_011000001001 : VALUE=19'b0000000_100010110101;
      15'b011_011000001010 : VALUE=19'b0000000_100010110101;
      15'b011_011000001011 : VALUE=19'b0000000_100010110101;
      15'b011_011000001100 : VALUE=19'b0000000_100010110101;
      15'b011_011000001101 : VALUE=19'b0000000_100010110101;
      15'b011_011000001110 : VALUE=19'b0000000_100010110100;
      15'b011_011000001111 : VALUE=19'b0000000_100010110100;
      15'b011_011000010000 : VALUE=19'b0000000_100010110100;
      15'b011_011000010001 : VALUE=19'b0000000_100010110100;
      15'b011_011000010010 : VALUE=19'b0000000_100010110100;
      15'b011_011000010011 : VALUE=19'b0000000_100010110100;
      15'b011_011000010100 : VALUE=19'b0000000_100010110100;
      15'b011_011000010101 : VALUE=19'b0000000_100010110100;
      15'b011_011000010110 : VALUE=19'b0000000_100010110100;
      15'b011_011000010111 : VALUE=19'b0000000_100010110100;
      15'b011_011000011000 : VALUE=19'b0000000_100010110100;
      15'b011_011000011001 : VALUE=19'b0000000_100010110100;
      15'b011_011000011010 : VALUE=19'b0000000_100010110011;
      15'b011_011000011011 : VALUE=19'b0000000_100010110011;
      15'b011_011000011100 : VALUE=19'b0000000_100010110011;
      15'b011_011000011101 : VALUE=19'b0000000_100010110011;
      15'b011_011000011110 : VALUE=19'b0000000_100010110011;
      15'b011_011000011111 : VALUE=19'b0000000_100010110011;
      15'b011_011000100000 : VALUE=19'b0000000_100010110011;
      15'b011_011000100001 : VALUE=19'b0000000_100010110011;
      15'b011_011000100010 : VALUE=19'b0000000_100010110011;
      15'b011_011000100011 : VALUE=19'b0000000_100010110011;
      15'b011_011000100100 : VALUE=19'b0000000_100010110011;
      15'b011_011000100101 : VALUE=19'b0000000_100010110011;
      15'b011_011000100110 : VALUE=19'b0000000_100010110011;
      15'b011_011000100111 : VALUE=19'b0000000_100010110010;
      15'b011_011000101000 : VALUE=19'b0000000_100010110010;
      15'b011_011000101001 : VALUE=19'b0000000_100010110010;
      15'b011_011000101010 : VALUE=19'b0000000_100010110010;
      15'b011_011000101011 : VALUE=19'b0000000_100010110010;
      15'b011_011000101100 : VALUE=19'b0000000_100010110010;
      15'b011_011000101101 : VALUE=19'b0000000_100010110010;
      15'b011_011000101110 : VALUE=19'b0000000_100010110010;
      15'b011_011000101111 : VALUE=19'b0000000_100010110010;
      15'b011_011000110000 : VALUE=19'b0000000_100010110010;
      15'b011_011000110001 : VALUE=19'b0000000_100010110010;
      15'b011_011000110010 : VALUE=19'b0000000_100010110010;
      15'b011_011000110011 : VALUE=19'b0000000_100010110001;
      15'b011_011000110100 : VALUE=19'b0000000_100010110001;
      15'b011_011000110101 : VALUE=19'b0000000_100010110001;
      15'b011_011000110110 : VALUE=19'b0000000_100010110001;
      15'b011_011000110111 : VALUE=19'b0000000_100010110001;
      15'b011_011000111000 : VALUE=19'b0000000_100010110001;
      15'b011_011000111001 : VALUE=19'b0000000_100010110001;
      15'b011_011000111010 : VALUE=19'b0000000_100010110001;
      15'b011_011000111011 : VALUE=19'b0000000_100010110001;
      15'b011_011000111100 : VALUE=19'b0000000_100010110001;
      15'b011_011000111101 : VALUE=19'b0000000_100010110001;
      15'b011_011000111110 : VALUE=19'b0000000_100010110001;
      15'b011_011000111111 : VALUE=19'b0000000_100010110001;
      15'b011_011001000000 : VALUE=19'b0000000_100010110000;
      15'b011_011001000001 : VALUE=19'b0000000_100010110000;
      15'b011_011001000010 : VALUE=19'b0000000_100010110000;
      15'b011_011001000011 : VALUE=19'b0000000_100010110000;
      15'b011_011001000100 : VALUE=19'b0000000_100010110000;
      15'b011_011001000101 : VALUE=19'b0000000_100010110000;
      15'b011_011001000110 : VALUE=19'b0000000_100010110000;
      15'b011_011001000111 : VALUE=19'b0000000_100010110000;
      15'b011_011001001000 : VALUE=19'b0000000_100010110000;
      15'b011_011001001001 : VALUE=19'b0000000_100010110000;
      15'b011_011001001010 : VALUE=19'b0000000_100010110000;
      15'b011_011001001011 : VALUE=19'b0000000_100010110000;
      15'b011_011001001100 : VALUE=19'b0000000_100010101111;
      15'b011_011001001101 : VALUE=19'b0000000_100010101111;
      15'b011_011001001110 : VALUE=19'b0000000_100010101111;
      15'b011_011001001111 : VALUE=19'b0000000_100010101111;
      15'b011_011001010000 : VALUE=19'b0000000_100010101111;
      15'b011_011001010001 : VALUE=19'b0000000_100010101111;
      15'b011_011001010010 : VALUE=19'b0000000_100010101111;
      15'b011_011001010011 : VALUE=19'b0000000_100010101111;
      15'b011_011001010100 : VALUE=19'b0000000_100010101111;
      15'b011_011001010101 : VALUE=19'b0000000_100010101111;
      15'b011_011001010110 : VALUE=19'b0000000_100010101111;
      15'b011_011001010111 : VALUE=19'b0000000_100010101111;
      15'b011_011001011000 : VALUE=19'b0000000_100010101111;
      15'b011_011001011001 : VALUE=19'b0000000_100010101110;
      15'b011_011001011010 : VALUE=19'b0000000_100010101110;
      15'b011_011001011011 : VALUE=19'b0000000_100010101110;
      15'b011_011001011100 : VALUE=19'b0000000_100010101110;
      15'b011_011001011101 : VALUE=19'b0000000_100010101110;
      15'b011_011001011110 : VALUE=19'b0000000_100010101110;
      15'b011_011001011111 : VALUE=19'b0000000_100010101110;
      15'b011_011001100000 : VALUE=19'b0000000_100010101110;
      15'b011_011001100001 : VALUE=19'b0000000_100010101110;
      15'b011_011001100010 : VALUE=19'b0000000_100010101110;
      15'b011_011001100011 : VALUE=19'b0000000_100010101110;
      15'b011_011001100100 : VALUE=19'b0000000_100010101110;
      15'b011_011001100101 : VALUE=19'b0000000_100010101101;
      15'b011_011001100110 : VALUE=19'b0000000_100010101101;
      15'b011_011001100111 : VALUE=19'b0000000_100010101101;
      15'b011_011001101000 : VALUE=19'b0000000_100010101101;
      15'b011_011001101001 : VALUE=19'b0000000_100010101101;
      15'b011_011001101010 : VALUE=19'b0000000_100010101101;
      15'b011_011001101011 : VALUE=19'b0000000_100010101101;
      15'b011_011001101100 : VALUE=19'b0000000_100010101101;
      15'b011_011001101101 : VALUE=19'b0000000_100010101101;
      15'b011_011001101110 : VALUE=19'b0000000_100010101101;
      15'b011_011001101111 : VALUE=19'b0000000_100010101101;
      15'b011_011001110000 : VALUE=19'b0000000_100010101101;
      15'b011_011001110001 : VALUE=19'b0000000_100010101101;
      15'b011_011001110010 : VALUE=19'b0000000_100010101100;
      15'b011_011001110011 : VALUE=19'b0000000_100010101100;
      15'b011_011001110100 : VALUE=19'b0000000_100010101100;
      15'b011_011001110101 : VALUE=19'b0000000_100010101100;
      15'b011_011001110110 : VALUE=19'b0000000_100010101100;
      15'b011_011001110111 : VALUE=19'b0000000_100010101100;
      15'b011_011001111000 : VALUE=19'b0000000_100010101100;
      15'b011_011001111001 : VALUE=19'b0000000_100010101100;
      15'b011_011001111010 : VALUE=19'b0000000_100010101100;
      15'b011_011001111011 : VALUE=19'b0000000_100010101100;
      15'b011_011001111100 : VALUE=19'b0000000_100010101100;
      15'b011_011001111101 : VALUE=19'b0000000_100010101100;
      15'b011_011001111110 : VALUE=19'b0000000_100010101011;
      15'b011_011001111111 : VALUE=19'b0000000_100010101011;
      15'b011_011010000000 : VALUE=19'b0000000_100010101011;
      15'b011_011010000001 : VALUE=19'b0000000_100010101011;
      15'b011_011010000010 : VALUE=19'b0000000_100010101011;
      15'b011_011010000011 : VALUE=19'b0000000_100010101011;
      15'b011_011010000100 : VALUE=19'b0000000_100010101011;
      15'b011_011010000101 : VALUE=19'b0000000_100010101011;
      15'b011_011010000110 : VALUE=19'b0000000_100010101011;
      15'b011_011010000111 : VALUE=19'b0000000_100010101011;
      15'b011_011010001000 : VALUE=19'b0000000_100010101011;
      15'b011_011010001001 : VALUE=19'b0000000_100010101011;
      15'b011_011010001010 : VALUE=19'b0000000_100010101011;
      15'b011_011010001011 : VALUE=19'b0000000_100010101010;
      15'b011_011010001100 : VALUE=19'b0000000_100010101010;
      15'b011_011010001101 : VALUE=19'b0000000_100010101010;
      15'b011_011010001110 : VALUE=19'b0000000_100010101010;
      15'b011_011010001111 : VALUE=19'b0000000_100010101010;
      15'b011_011010010000 : VALUE=19'b0000000_100010101010;
      15'b011_011010010001 : VALUE=19'b0000000_100010101010;
      15'b011_011010010010 : VALUE=19'b0000000_100010101010;
      15'b011_011010010011 : VALUE=19'b0000000_100010101010;
      15'b011_011010010100 : VALUE=19'b0000000_100010101010;
      15'b011_011010010101 : VALUE=19'b0000000_100010101010;
      15'b011_011010010110 : VALUE=19'b0000000_100010101010;
      15'b011_011010010111 : VALUE=19'b0000000_100010101010;
      15'b011_011010011000 : VALUE=19'b0000000_100010101001;
      15'b011_011010011001 : VALUE=19'b0000000_100010101001;
      15'b011_011010011010 : VALUE=19'b0000000_100010101001;
      15'b011_011010011011 : VALUE=19'b0000000_100010101001;
      15'b011_011010011100 : VALUE=19'b0000000_100010101001;
      15'b011_011010011101 : VALUE=19'b0000000_100010101001;
      15'b011_011010011110 : VALUE=19'b0000000_100010101001;
      15'b011_011010011111 : VALUE=19'b0000000_100010101001;
      15'b011_011010100000 : VALUE=19'b0000000_100010101001;
      15'b011_011010100001 : VALUE=19'b0000000_100010101001;
      15'b011_011010100010 : VALUE=19'b0000000_100010101001;
      15'b011_011010100011 : VALUE=19'b0000000_100010101001;
      15'b011_011010100100 : VALUE=19'b0000000_100010101000;
      15'b011_011010100101 : VALUE=19'b0000000_100010101000;
      15'b011_011010100110 : VALUE=19'b0000000_100010101000;
      15'b011_011010100111 : VALUE=19'b0000000_100010101000;
      15'b011_011010101000 : VALUE=19'b0000000_100010101000;
      15'b011_011010101001 : VALUE=19'b0000000_100010101000;
      15'b011_011010101010 : VALUE=19'b0000000_100010101000;
      15'b011_011010101011 : VALUE=19'b0000000_100010101000;
      15'b011_011010101100 : VALUE=19'b0000000_100010101000;
      15'b011_011010101101 : VALUE=19'b0000000_100010101000;
      15'b011_011010101110 : VALUE=19'b0000000_100010101000;
      15'b011_011010101111 : VALUE=19'b0000000_100010101000;
      15'b011_011010110000 : VALUE=19'b0000000_100010101000;
      15'b011_011010110001 : VALUE=19'b0000000_100010100111;
      15'b011_011010110010 : VALUE=19'b0000000_100010100111;
      15'b011_011010110011 : VALUE=19'b0000000_100010100111;
      15'b011_011010110100 : VALUE=19'b0000000_100010100111;
      15'b011_011010110101 : VALUE=19'b0000000_100010100111;
      15'b011_011010110110 : VALUE=19'b0000000_100010100111;
      15'b011_011010110111 : VALUE=19'b0000000_100010100111;
      15'b011_011010111000 : VALUE=19'b0000000_100010100111;
      15'b011_011010111001 : VALUE=19'b0000000_100010100111;
      15'b011_011010111010 : VALUE=19'b0000000_100010100111;
      15'b011_011010111011 : VALUE=19'b0000000_100010100111;
      15'b011_011010111100 : VALUE=19'b0000000_100010100111;
      15'b011_011010111101 : VALUE=19'b0000000_100010100110;
      15'b011_011010111110 : VALUE=19'b0000000_100010100110;
      15'b011_011010111111 : VALUE=19'b0000000_100010100110;
      15'b011_011011000000 : VALUE=19'b0000000_100010100110;
      15'b011_011011000001 : VALUE=19'b0000000_100010100110;
      15'b011_011011000010 : VALUE=19'b0000000_100010100110;
      15'b011_011011000011 : VALUE=19'b0000000_100010100110;
      15'b011_011011000100 : VALUE=19'b0000000_100010100110;
      15'b011_011011000101 : VALUE=19'b0000000_100010100110;
      15'b011_011011000110 : VALUE=19'b0000000_100010100110;
      15'b011_011011000111 : VALUE=19'b0000000_100010100110;
      15'b011_011011001000 : VALUE=19'b0000000_100010100110;
      15'b011_011011001001 : VALUE=19'b0000000_100010100110;
      15'b011_011011001010 : VALUE=19'b0000000_100010100101;
      15'b011_011011001011 : VALUE=19'b0000000_100010100101;
      15'b011_011011001100 : VALUE=19'b0000000_100010100101;
      15'b011_011011001101 : VALUE=19'b0000000_100010100101;
      15'b011_011011001110 : VALUE=19'b0000000_100010100101;
      15'b011_011011001111 : VALUE=19'b0000000_100010100101;
      15'b011_011011010000 : VALUE=19'b0000000_100010100101;
      15'b011_011011010001 : VALUE=19'b0000000_100010100101;
      15'b011_011011010010 : VALUE=19'b0000000_100010100101;
      15'b011_011011010011 : VALUE=19'b0000000_100010100101;
      15'b011_011011010100 : VALUE=19'b0000000_100010100101;
      15'b011_011011010101 : VALUE=19'b0000000_100010100101;
      15'b011_011011010110 : VALUE=19'b0000000_100010100101;
      15'b011_011011010111 : VALUE=19'b0000000_100010100100;
      15'b011_011011011000 : VALUE=19'b0000000_100010100100;
      15'b011_011011011001 : VALUE=19'b0000000_100010100100;
      15'b011_011011011010 : VALUE=19'b0000000_100010100100;
      15'b011_011011011011 : VALUE=19'b0000000_100010100100;
      15'b011_011011011100 : VALUE=19'b0000000_100010100100;
      15'b011_011011011101 : VALUE=19'b0000000_100010100100;
      15'b011_011011011110 : VALUE=19'b0000000_100010100100;
      15'b011_011011011111 : VALUE=19'b0000000_100010100100;
      15'b011_011011100000 : VALUE=19'b0000000_100010100100;
      15'b011_011011100001 : VALUE=19'b0000000_100010100100;
      15'b011_011011100010 : VALUE=19'b0000000_100010100100;
      15'b011_011011100011 : VALUE=19'b0000000_100010100011;
      15'b011_011011100100 : VALUE=19'b0000000_100010100011;
      15'b011_011011100101 : VALUE=19'b0000000_100010100011;
      15'b011_011011100110 : VALUE=19'b0000000_100010100011;
      15'b011_011011100111 : VALUE=19'b0000000_100010100011;
      15'b011_011011101000 : VALUE=19'b0000000_100010100011;
      15'b011_011011101001 : VALUE=19'b0000000_100010100011;
      15'b011_011011101010 : VALUE=19'b0000000_100010100011;
      15'b011_011011101011 : VALUE=19'b0000000_100010100011;
      15'b011_011011101100 : VALUE=19'b0000000_100010100011;
      15'b011_011011101101 : VALUE=19'b0000000_100010100011;
      15'b011_011011101110 : VALUE=19'b0000000_100010100011;
      15'b011_011011101111 : VALUE=19'b0000000_100010100011;
      15'b011_011011110000 : VALUE=19'b0000000_100010100010;
      15'b011_011011110001 : VALUE=19'b0000000_100010100010;
      15'b011_011011110010 : VALUE=19'b0000000_100010100010;
      15'b011_011011110011 : VALUE=19'b0000000_100010100010;
      15'b011_011011110100 : VALUE=19'b0000000_100010100010;
      15'b011_011011110101 : VALUE=19'b0000000_100010100010;
      15'b011_011011110110 : VALUE=19'b0000000_100010100010;
      15'b011_011011110111 : VALUE=19'b0000000_100010100010;
      15'b011_011011111000 : VALUE=19'b0000000_100010100010;
      15'b011_011011111001 : VALUE=19'b0000000_100010100010;
      15'b011_011011111010 : VALUE=19'b0000000_100010100010;
      15'b011_011011111011 : VALUE=19'b0000000_100010100010;
      15'b011_011011111100 : VALUE=19'b0000000_100010100010;
      15'b011_011011111101 : VALUE=19'b0000000_100010100001;
      15'b011_011011111110 : VALUE=19'b0000000_100010100001;
      15'b011_011011111111 : VALUE=19'b0000000_100010100001;
      15'b011_011100000000 : VALUE=19'b0000000_100010100001;
      15'b011_011100000001 : VALUE=19'b0000000_100010100001;
      15'b011_011100000010 : VALUE=19'b0000000_100010100001;
      15'b011_011100000011 : VALUE=19'b0000000_100010100001;
      15'b011_011100000100 : VALUE=19'b0000000_100010100001;
      15'b011_011100000101 : VALUE=19'b0000000_100010100001;
      15'b011_011100000110 : VALUE=19'b0000000_100010100001;
      15'b011_011100000111 : VALUE=19'b0000000_100010100001;
      15'b011_011100001000 : VALUE=19'b0000000_100010100001;
      15'b011_011100001001 : VALUE=19'b0000000_100010100001;
      15'b011_011100001010 : VALUE=19'b0000000_100010100000;
      15'b011_011100001011 : VALUE=19'b0000000_100010100000;
      15'b011_011100001100 : VALUE=19'b0000000_100010100000;
      15'b011_011100001101 : VALUE=19'b0000000_100010100000;
      15'b011_011100001110 : VALUE=19'b0000000_100010100000;
      15'b011_011100001111 : VALUE=19'b0000000_100010100000;
      15'b011_011100010000 : VALUE=19'b0000000_100010100000;
      15'b011_011100010001 : VALUE=19'b0000000_100010100000;
      15'b011_011100010010 : VALUE=19'b0000000_100010100000;
      15'b011_011100010011 : VALUE=19'b0000000_100010100000;
      15'b011_011100010100 : VALUE=19'b0000000_100010100000;
      15'b011_011100010101 : VALUE=19'b0000000_100010100000;
      15'b011_011100010110 : VALUE=19'b0000000_100010011111;
      15'b011_011100010111 : VALUE=19'b0000000_100010011111;
      15'b011_011100011000 : VALUE=19'b0000000_100010011111;
      15'b011_011100011001 : VALUE=19'b0000000_100010011111;
      15'b011_011100011010 : VALUE=19'b0000000_100010011111;
      15'b011_011100011011 : VALUE=19'b0000000_100010011111;
      15'b011_011100011100 : VALUE=19'b0000000_100010011111;
      15'b011_011100011101 : VALUE=19'b0000000_100010011111;
      15'b011_011100011110 : VALUE=19'b0000000_100010011111;
      15'b011_011100011111 : VALUE=19'b0000000_100010011111;
      15'b011_011100100000 : VALUE=19'b0000000_100010011111;
      15'b011_011100100001 : VALUE=19'b0000000_100010011111;
      15'b011_011100100010 : VALUE=19'b0000000_100010011111;
      15'b011_011100100011 : VALUE=19'b0000000_100010011110;
      15'b011_011100100100 : VALUE=19'b0000000_100010011110;
      15'b011_011100100101 : VALUE=19'b0000000_100010011110;
      15'b011_011100100110 : VALUE=19'b0000000_100010011110;
      15'b011_011100100111 : VALUE=19'b0000000_100010011110;
      15'b011_011100101000 : VALUE=19'b0000000_100010011110;
      15'b011_011100101001 : VALUE=19'b0000000_100010011110;
      15'b011_011100101010 : VALUE=19'b0000000_100010011110;
      15'b011_011100101011 : VALUE=19'b0000000_100010011110;
      15'b011_011100101100 : VALUE=19'b0000000_100010011110;
      15'b011_011100101101 : VALUE=19'b0000000_100010011110;
      15'b011_011100101110 : VALUE=19'b0000000_100010011110;
      15'b011_011100101111 : VALUE=19'b0000000_100010011110;
      15'b011_011100110000 : VALUE=19'b0000000_100010011101;
      15'b011_011100110001 : VALUE=19'b0000000_100010011101;
      15'b011_011100110010 : VALUE=19'b0000000_100010011101;
      15'b011_011100110011 : VALUE=19'b0000000_100010011101;
      15'b011_011100110100 : VALUE=19'b0000000_100010011101;
      15'b011_011100110101 : VALUE=19'b0000000_100010011101;
      15'b011_011100110110 : VALUE=19'b0000000_100010011101;
      15'b011_011100110111 : VALUE=19'b0000000_100010011101;
      15'b011_011100111000 : VALUE=19'b0000000_100010011101;
      15'b011_011100111001 : VALUE=19'b0000000_100010011101;
      15'b011_011100111010 : VALUE=19'b0000000_100010011101;
      15'b011_011100111011 : VALUE=19'b0000000_100010011101;
      15'b011_011100111100 : VALUE=19'b0000000_100010011101;
      15'b011_011100111101 : VALUE=19'b0000000_100010011100;
      15'b011_011100111110 : VALUE=19'b0000000_100010011100;
      15'b011_011100111111 : VALUE=19'b0000000_100010011100;
      15'b011_011101000000 : VALUE=19'b0000000_100010011100;
      15'b011_011101000001 : VALUE=19'b0000000_100010011100;
      15'b011_011101000010 : VALUE=19'b0000000_100010011100;
      15'b011_011101000011 : VALUE=19'b0000000_100010011100;
      15'b011_011101000100 : VALUE=19'b0000000_100010011100;
      15'b011_011101000101 : VALUE=19'b0000000_100010011100;
      15'b011_011101000110 : VALUE=19'b0000000_100010011100;
      15'b011_011101000111 : VALUE=19'b0000000_100010011100;
      15'b011_011101001000 : VALUE=19'b0000000_100010011100;
      15'b011_011101001001 : VALUE=19'b0000000_100010011100;
      15'b011_011101001010 : VALUE=19'b0000000_100010011011;
      15'b011_011101001011 : VALUE=19'b0000000_100010011011;
      15'b011_011101001100 : VALUE=19'b0000000_100010011011;
      15'b011_011101001101 : VALUE=19'b0000000_100010011011;
      15'b011_011101001110 : VALUE=19'b0000000_100010011011;
      15'b011_011101001111 : VALUE=19'b0000000_100010011011;
      15'b011_011101010000 : VALUE=19'b0000000_100010011011;
      15'b011_011101010001 : VALUE=19'b0000000_100010011011;
      15'b011_011101010010 : VALUE=19'b0000000_100010011011;
      15'b011_011101010011 : VALUE=19'b0000000_100010011011;
      15'b011_011101010100 : VALUE=19'b0000000_100010011011;
      15'b011_011101010101 : VALUE=19'b0000000_100010011011;
      15'b011_011101010110 : VALUE=19'b0000000_100010011011;
      15'b011_011101010111 : VALUE=19'b0000000_100010011010;
      15'b011_011101011000 : VALUE=19'b0000000_100010011010;
      15'b011_011101011001 : VALUE=19'b0000000_100010011010;
      15'b011_011101011010 : VALUE=19'b0000000_100010011010;
      15'b011_011101011011 : VALUE=19'b0000000_100010011010;
      15'b011_011101011100 : VALUE=19'b0000000_100010011010;
      15'b011_011101011101 : VALUE=19'b0000000_100010011010;
      15'b011_011101011110 : VALUE=19'b0000000_100010011010;
      15'b011_011101011111 : VALUE=19'b0000000_100010011010;
      15'b011_011101100000 : VALUE=19'b0000000_100010011010;
      15'b011_011101100001 : VALUE=19'b0000000_100010011010;
      15'b011_011101100010 : VALUE=19'b0000000_100010011010;
      15'b011_011101100011 : VALUE=19'b0000000_100010011001;
      15'b011_011101100100 : VALUE=19'b0000000_100010011001;
      15'b011_011101100101 : VALUE=19'b0000000_100010011001;
      15'b011_011101100110 : VALUE=19'b0000000_100010011001;
      15'b011_011101100111 : VALUE=19'b0000000_100010011001;
      15'b011_011101101000 : VALUE=19'b0000000_100010011001;
      15'b011_011101101001 : VALUE=19'b0000000_100010011001;
      15'b011_011101101010 : VALUE=19'b0000000_100010011001;
      15'b011_011101101011 : VALUE=19'b0000000_100010011001;
      15'b011_011101101100 : VALUE=19'b0000000_100010011001;
      15'b011_011101101101 : VALUE=19'b0000000_100010011001;
      15'b011_011101101110 : VALUE=19'b0000000_100010011001;
      15'b011_011101101111 : VALUE=19'b0000000_100010011001;
      15'b011_011101110000 : VALUE=19'b0000000_100010011000;
      15'b011_011101110001 : VALUE=19'b0000000_100010011000;
      15'b011_011101110010 : VALUE=19'b0000000_100010011000;
      15'b011_011101110011 : VALUE=19'b0000000_100010011000;
      15'b011_011101110100 : VALUE=19'b0000000_100010011000;
      15'b011_011101110101 : VALUE=19'b0000000_100010011000;
      15'b011_011101110110 : VALUE=19'b0000000_100010011000;
      15'b011_011101110111 : VALUE=19'b0000000_100010011000;
      15'b011_011101111000 : VALUE=19'b0000000_100010011000;
      15'b011_011101111001 : VALUE=19'b0000000_100010011000;
      15'b011_011101111010 : VALUE=19'b0000000_100010011000;
      15'b011_011101111011 : VALUE=19'b0000000_100010011000;
      15'b011_011101111100 : VALUE=19'b0000000_100010011000;
      15'b011_011101111101 : VALUE=19'b0000000_100010010111;
      15'b011_011101111110 : VALUE=19'b0000000_100010010111;
      15'b011_011101111111 : VALUE=19'b0000000_100010010111;
      15'b011_011110000000 : VALUE=19'b0000000_100010010111;
      15'b011_011110000001 : VALUE=19'b0000000_100010010111;
      15'b011_011110000010 : VALUE=19'b0000000_100010010111;
      15'b011_011110000011 : VALUE=19'b0000000_100010010111;
      15'b011_011110000100 : VALUE=19'b0000000_100010010111;
      15'b011_011110000101 : VALUE=19'b0000000_100010010111;
      15'b011_011110000110 : VALUE=19'b0000000_100010010111;
      15'b011_011110000111 : VALUE=19'b0000000_100010010111;
      15'b011_011110001000 : VALUE=19'b0000000_100010010111;
      15'b011_011110001001 : VALUE=19'b0000000_100010010111;
      15'b011_011110001010 : VALUE=19'b0000000_100010010110;
      15'b011_011110001011 : VALUE=19'b0000000_100010010110;
      15'b011_011110001100 : VALUE=19'b0000000_100010010110;
      15'b011_011110001101 : VALUE=19'b0000000_100010010110;
      15'b011_011110001110 : VALUE=19'b0000000_100010010110;
      15'b011_011110001111 : VALUE=19'b0000000_100010010110;
      15'b011_011110010000 : VALUE=19'b0000000_100010010110;
      15'b011_011110010001 : VALUE=19'b0000000_100010010110;
      15'b011_011110010010 : VALUE=19'b0000000_100010010110;
      15'b011_011110010011 : VALUE=19'b0000000_100010010110;
      15'b011_011110010100 : VALUE=19'b0000000_100010010110;
      15'b011_011110010101 : VALUE=19'b0000000_100010010110;
      15'b011_011110010110 : VALUE=19'b0000000_100010010110;
      15'b011_011110010111 : VALUE=19'b0000000_100010010101;
      15'b011_011110011000 : VALUE=19'b0000000_100010010101;
      15'b011_011110011001 : VALUE=19'b0000000_100010010101;
      15'b011_011110011010 : VALUE=19'b0000000_100010010101;
      15'b011_011110011011 : VALUE=19'b0000000_100010010101;
      15'b011_011110011100 : VALUE=19'b0000000_100010010101;
      15'b011_011110011101 : VALUE=19'b0000000_100010010101;
      15'b011_011110011110 : VALUE=19'b0000000_100010010101;
      15'b011_011110011111 : VALUE=19'b0000000_100010010101;
      15'b011_011110100000 : VALUE=19'b0000000_100010010101;
      15'b011_011110100001 : VALUE=19'b0000000_100010010101;
      15'b011_011110100010 : VALUE=19'b0000000_100010010101;
      15'b011_011110100011 : VALUE=19'b0000000_100010010101;
      15'b011_011110100100 : VALUE=19'b0000000_100010010100;
      15'b011_011110100101 : VALUE=19'b0000000_100010010100;
      15'b011_011110100110 : VALUE=19'b0000000_100010010100;
      15'b011_011110100111 : VALUE=19'b0000000_100010010100;
      15'b011_011110101000 : VALUE=19'b0000000_100010010100;
      15'b011_011110101001 : VALUE=19'b0000000_100010010100;
      15'b011_011110101010 : VALUE=19'b0000000_100010010100;
      15'b011_011110101011 : VALUE=19'b0000000_100010010100;
      15'b011_011110101100 : VALUE=19'b0000000_100010010100;
      15'b011_011110101101 : VALUE=19'b0000000_100010010100;
      15'b011_011110101110 : VALUE=19'b0000000_100010010100;
      15'b011_011110101111 : VALUE=19'b0000000_100010010100;
      15'b011_011110110000 : VALUE=19'b0000000_100010010100;
      15'b011_011110110001 : VALUE=19'b0000000_100010010011;
      15'b011_011110110010 : VALUE=19'b0000000_100010010011;
      15'b011_011110110011 : VALUE=19'b0000000_100010010011;
      15'b011_011110110100 : VALUE=19'b0000000_100010010011;
      15'b011_011110110101 : VALUE=19'b0000000_100010010011;
      15'b011_011110110110 : VALUE=19'b0000000_100010010011;
      15'b011_011110110111 : VALUE=19'b0000000_100010010011;
      15'b011_011110111000 : VALUE=19'b0000000_100010010011;
      15'b011_011110111001 : VALUE=19'b0000000_100010010011;
      15'b011_011110111010 : VALUE=19'b0000000_100010010011;
      15'b011_011110111011 : VALUE=19'b0000000_100010010011;
      15'b011_011110111100 : VALUE=19'b0000000_100010010011;
      15'b011_011110111101 : VALUE=19'b0000000_100010010011;
      15'b011_011110111110 : VALUE=19'b0000000_100010010010;
      15'b011_011110111111 : VALUE=19'b0000000_100010010010;
      15'b011_011111000000 : VALUE=19'b0000000_100010010010;
      15'b011_011111000001 : VALUE=19'b0000000_100010010010;
      15'b011_011111000010 : VALUE=19'b0000000_100010010010;
      15'b011_011111000011 : VALUE=19'b0000000_100010010010;
      15'b011_011111000100 : VALUE=19'b0000000_100010010010;
      15'b011_011111000101 : VALUE=19'b0000000_100010010010;
      15'b011_011111000110 : VALUE=19'b0000000_100010010010;
      15'b011_011111000111 : VALUE=19'b0000000_100010010010;
      15'b011_011111001000 : VALUE=19'b0000000_100010010010;
      15'b011_011111001001 : VALUE=19'b0000000_100010010010;
      15'b011_011111001010 : VALUE=19'b0000000_100010010010;
      15'b011_011111001011 : VALUE=19'b0000000_100010010001;
      15'b011_011111001100 : VALUE=19'b0000000_100010010001;
      15'b011_011111001101 : VALUE=19'b0000000_100010010001;
      15'b011_011111001110 : VALUE=19'b0000000_100010010001;
      15'b011_011111001111 : VALUE=19'b0000000_100010010001;
      15'b011_011111010000 : VALUE=19'b0000000_100010010001;
      15'b011_011111010001 : VALUE=19'b0000000_100010010001;
      15'b011_011111010010 : VALUE=19'b0000000_100010010001;
      15'b011_011111010011 : VALUE=19'b0000000_100010010001;
      15'b011_011111010100 : VALUE=19'b0000000_100010010001;
      15'b011_011111010101 : VALUE=19'b0000000_100010010001;
      15'b011_011111010110 : VALUE=19'b0000000_100010010001;
      15'b011_011111010111 : VALUE=19'b0000000_100010010001;
      15'b011_011111011000 : VALUE=19'b0000000_100010010000;
      15'b011_011111011001 : VALUE=19'b0000000_100010010000;
      15'b011_011111011010 : VALUE=19'b0000000_100010010000;
      15'b011_011111011011 : VALUE=19'b0000000_100010010000;
      15'b011_011111011100 : VALUE=19'b0000000_100010010000;
      15'b011_011111011101 : VALUE=19'b0000000_100010010000;
      15'b011_011111011110 : VALUE=19'b0000000_100010010000;
      15'b011_011111011111 : VALUE=19'b0000000_100010010000;
      15'b011_011111100000 : VALUE=19'b0000000_100010010000;
      15'b011_011111100001 : VALUE=19'b0000000_100010010000;
      15'b011_011111100010 : VALUE=19'b0000000_100010010000;
      15'b011_011111100011 : VALUE=19'b0000000_100010010000;
      15'b011_011111100100 : VALUE=19'b0000000_100010010000;
      15'b011_011111100101 : VALUE=19'b0000000_100010001111;
      15'b011_011111100110 : VALUE=19'b0000000_100010001111;
      15'b011_011111100111 : VALUE=19'b0000000_100010001111;
      15'b011_011111101000 : VALUE=19'b0000000_100010001111;
      15'b011_011111101001 : VALUE=19'b0000000_100010001111;
      15'b011_011111101010 : VALUE=19'b0000000_100010001111;
      15'b011_011111101011 : VALUE=19'b0000000_100010001111;
      15'b011_011111101100 : VALUE=19'b0000000_100010001111;
      15'b011_011111101101 : VALUE=19'b0000000_100010001111;
      15'b011_011111101110 : VALUE=19'b0000000_100010001111;
      15'b011_011111101111 : VALUE=19'b0000000_100010001111;
      15'b011_011111110000 : VALUE=19'b0000000_100010001111;
      15'b011_011111110001 : VALUE=19'b0000000_100010001111;
      15'b011_011111110010 : VALUE=19'b0000000_100010001110;
      15'b011_011111110011 : VALUE=19'b0000000_100010001110;
      15'b011_011111110100 : VALUE=19'b0000000_100010001110;
      15'b011_011111110101 : VALUE=19'b0000000_100010001110;
      15'b011_011111110110 : VALUE=19'b0000000_100010001110;
      15'b011_011111110111 : VALUE=19'b0000000_100010001110;
      15'b011_011111111000 : VALUE=19'b0000000_100010001110;
      15'b011_011111111001 : VALUE=19'b0000000_100010001110;
      15'b011_011111111010 : VALUE=19'b0000000_100010001110;
      15'b011_011111111011 : VALUE=19'b0000000_100010001110;
      15'b011_011111111100 : VALUE=19'b0000000_100010001110;
      15'b011_011111111101 : VALUE=19'b0000000_100010001110;
      15'b011_011111111110 : VALUE=19'b0000000_100010001110;
      15'b011_011111111111 : VALUE=19'b0000000_100010001101;
      15'b011_100000000000 : VALUE=19'b0000000_100010001101;
      15'b011_100000000001 : VALUE=19'b0000000_100010001101;
      15'b011_100000000010 : VALUE=19'b0000000_100010001101;
      15'b011_100000000011 : VALUE=19'b0000000_100010001101;
      15'b011_100000000100 : VALUE=19'b0000000_100010001101;
      15'b011_100000000101 : VALUE=19'b0000000_100010001101;
      15'b011_100000000110 : VALUE=19'b0000000_100010001101;
      15'b011_100000000111 : VALUE=19'b0000000_100010001101;
      15'b011_100000001000 : VALUE=19'b0000000_100010001101;
      15'b011_100000001001 : VALUE=19'b0000000_100010001101;
      15'b011_100000001010 : VALUE=19'b0000000_100010001101;
      15'b011_100000001011 : VALUE=19'b0000000_100010001101;
      15'b011_100000001100 : VALUE=19'b0000000_100010001100;
      15'b011_100000001101 : VALUE=19'b0000000_100010001100;
      15'b011_100000001110 : VALUE=19'b0000000_100010001100;
      15'b011_100000001111 : VALUE=19'b0000000_100010001100;
      15'b011_100000010000 : VALUE=19'b0000000_100010001100;
      15'b011_100000010001 : VALUE=19'b0000000_100010001100;
      15'b011_100000010010 : VALUE=19'b0000000_100010001100;
      15'b011_100000010011 : VALUE=19'b0000000_100010001100;
      15'b011_100000010100 : VALUE=19'b0000000_100010001100;
      15'b011_100000010101 : VALUE=19'b0000000_100010001100;
      15'b011_100000010110 : VALUE=19'b0000000_100010001100;
      15'b011_100000010111 : VALUE=19'b0000000_100010001100;
      15'b011_100000011000 : VALUE=19'b0000000_100010001100;
      15'b011_100000011001 : VALUE=19'b0000000_100010001011;
      15'b011_100000011010 : VALUE=19'b0000000_100010001011;
      15'b011_100000011011 : VALUE=19'b0000000_100010001011;
      15'b011_100000011100 : VALUE=19'b0000000_100010001011;
      15'b011_100000011101 : VALUE=19'b0000000_100010001011;
      15'b011_100000011110 : VALUE=19'b0000000_100010001011;
      15'b011_100000011111 : VALUE=19'b0000000_100010001011;
      15'b011_100000100000 : VALUE=19'b0000000_100010001011;
      15'b011_100000100001 : VALUE=19'b0000000_100010001011;
      15'b011_100000100010 : VALUE=19'b0000000_100010001011;
      15'b011_100000100011 : VALUE=19'b0000000_100010001011;
      15'b011_100000100100 : VALUE=19'b0000000_100010001011;
      15'b011_100000100101 : VALUE=19'b0000000_100010001011;
      15'b011_100000100110 : VALUE=19'b0000000_100010001011;
      15'b011_100000100111 : VALUE=19'b0000000_100010001010;
      15'b011_100000101000 : VALUE=19'b0000000_100010001010;
      15'b011_100000101001 : VALUE=19'b0000000_100010001010;
      15'b011_100000101010 : VALUE=19'b0000000_100010001010;
      15'b011_100000101011 : VALUE=19'b0000000_100010001010;
      15'b011_100000101100 : VALUE=19'b0000000_100010001010;
      15'b011_100000101101 : VALUE=19'b0000000_100010001010;
      15'b011_100000101110 : VALUE=19'b0000000_100010001010;
      15'b011_100000101111 : VALUE=19'b0000000_100010001010;
      15'b011_100000110000 : VALUE=19'b0000000_100010001010;
      15'b011_100000110001 : VALUE=19'b0000000_100010001010;
      15'b011_100000110010 : VALUE=19'b0000000_100010001010;
      15'b011_100000110011 : VALUE=19'b0000000_100010001010;
      15'b011_100000110100 : VALUE=19'b0000000_100010001001;
      15'b011_100000110101 : VALUE=19'b0000000_100010001001;
      15'b011_100000110110 : VALUE=19'b0000000_100010001001;
      15'b011_100000110111 : VALUE=19'b0000000_100010001001;
      15'b011_100000111000 : VALUE=19'b0000000_100010001001;
      15'b011_100000111001 : VALUE=19'b0000000_100010001001;
      15'b011_100000111010 : VALUE=19'b0000000_100010001001;
      15'b011_100000111011 : VALUE=19'b0000000_100010001001;
      15'b011_100000111100 : VALUE=19'b0000000_100010001001;
      15'b011_100000111101 : VALUE=19'b0000000_100010001001;
      15'b011_100000111110 : VALUE=19'b0000000_100010001001;
      15'b011_100000111111 : VALUE=19'b0000000_100010001001;
      15'b011_100001000000 : VALUE=19'b0000000_100010001001;
      15'b011_100001000001 : VALUE=19'b0000000_100010001000;
      15'b011_100001000010 : VALUE=19'b0000000_100010001000;
      15'b011_100001000011 : VALUE=19'b0000000_100010001000;
      15'b011_100001000100 : VALUE=19'b0000000_100010001000;
      15'b011_100001000101 : VALUE=19'b0000000_100010001000;
      15'b011_100001000110 : VALUE=19'b0000000_100010001000;
      15'b011_100001000111 : VALUE=19'b0000000_100010001000;
      15'b011_100001001000 : VALUE=19'b0000000_100010001000;
      15'b011_100001001001 : VALUE=19'b0000000_100010001000;
      15'b011_100001001010 : VALUE=19'b0000000_100010001000;
      15'b011_100001001011 : VALUE=19'b0000000_100010001000;
      15'b011_100001001100 : VALUE=19'b0000000_100010001000;
      15'b011_100001001101 : VALUE=19'b0000000_100010001000;
      15'b011_100001001110 : VALUE=19'b0000000_100010000111;
      15'b011_100001001111 : VALUE=19'b0000000_100010000111;
      15'b011_100001010000 : VALUE=19'b0000000_100010000111;
      15'b011_100001010001 : VALUE=19'b0000000_100010000111;
      15'b011_100001010010 : VALUE=19'b0000000_100010000111;
      15'b011_100001010011 : VALUE=19'b0000000_100010000111;
      15'b011_100001010100 : VALUE=19'b0000000_100010000111;
      15'b011_100001010101 : VALUE=19'b0000000_100010000111;
      15'b011_100001010110 : VALUE=19'b0000000_100010000111;
      15'b011_100001010111 : VALUE=19'b0000000_100010000111;
      15'b011_100001011000 : VALUE=19'b0000000_100010000111;
      15'b011_100001011001 : VALUE=19'b0000000_100010000111;
      15'b011_100001011010 : VALUE=19'b0000000_100010000111;
      15'b011_100001011011 : VALUE=19'b0000000_100010000110;
      15'b011_100001011100 : VALUE=19'b0000000_100010000110;
      15'b011_100001011101 : VALUE=19'b0000000_100010000110;
      15'b011_100001011110 : VALUE=19'b0000000_100010000110;
      15'b011_100001011111 : VALUE=19'b0000000_100010000110;
      15'b011_100001100000 : VALUE=19'b0000000_100010000110;
      15'b011_100001100001 : VALUE=19'b0000000_100010000110;
      15'b011_100001100010 : VALUE=19'b0000000_100010000110;
      15'b011_100001100011 : VALUE=19'b0000000_100010000110;
      15'b011_100001100100 : VALUE=19'b0000000_100010000110;
      15'b011_100001100101 : VALUE=19'b0000000_100010000110;
      15'b011_100001100110 : VALUE=19'b0000000_100010000110;
      15'b011_100001100111 : VALUE=19'b0000000_100010000110;
      15'b011_100001101000 : VALUE=19'b0000000_100010000110;
      15'b011_100001101001 : VALUE=19'b0000000_100010000101;
      15'b011_100001101010 : VALUE=19'b0000000_100010000101;
      15'b011_100001101011 : VALUE=19'b0000000_100010000101;
      15'b011_100001101100 : VALUE=19'b0000000_100010000101;
      15'b011_100001101101 : VALUE=19'b0000000_100010000101;
      15'b011_100001101110 : VALUE=19'b0000000_100010000101;
      15'b011_100001101111 : VALUE=19'b0000000_100010000101;
      15'b011_100001110000 : VALUE=19'b0000000_100010000101;
      15'b011_100001110001 : VALUE=19'b0000000_100010000101;
      15'b011_100001110010 : VALUE=19'b0000000_100010000101;
      15'b011_100001110011 : VALUE=19'b0000000_100010000101;
      15'b011_100001110100 : VALUE=19'b0000000_100010000101;
      15'b011_100001110101 : VALUE=19'b0000000_100010000101;
      15'b011_100001110110 : VALUE=19'b0000000_100010000100;
      15'b011_100001110111 : VALUE=19'b0000000_100010000100;
      15'b011_100001111000 : VALUE=19'b0000000_100010000100;
      15'b011_100001111001 : VALUE=19'b0000000_100010000100;
      15'b011_100001111010 : VALUE=19'b0000000_100010000100;
      15'b011_100001111011 : VALUE=19'b0000000_100010000100;
      15'b011_100001111100 : VALUE=19'b0000000_100010000100;
      15'b011_100001111101 : VALUE=19'b0000000_100010000100;
      15'b011_100001111110 : VALUE=19'b0000000_100010000100;
      15'b011_100001111111 : VALUE=19'b0000000_100010000100;
      15'b011_100010000000 : VALUE=19'b0000000_100010000100;
      15'b011_100010000001 : VALUE=19'b0000000_100010000100;
      15'b011_100010000010 : VALUE=19'b0000000_100010000100;
      15'b011_100010000011 : VALUE=19'b0000000_100010000011;
      15'b011_100010000100 : VALUE=19'b0000000_100010000011;
      15'b011_100010000101 : VALUE=19'b0000000_100010000011;
      15'b011_100010000110 : VALUE=19'b0000000_100010000011;
      15'b011_100010000111 : VALUE=19'b0000000_100010000011;
      15'b011_100010001000 : VALUE=19'b0000000_100010000011;
      15'b011_100010001001 : VALUE=19'b0000000_100010000011;
      15'b011_100010001010 : VALUE=19'b0000000_100010000011;
      15'b011_100010001011 : VALUE=19'b0000000_100010000011;
      15'b011_100010001100 : VALUE=19'b0000000_100010000011;
      15'b011_100010001101 : VALUE=19'b0000000_100010000011;
      15'b011_100010001110 : VALUE=19'b0000000_100010000011;
      15'b011_100010001111 : VALUE=19'b0000000_100010000011;
      15'b011_100010010000 : VALUE=19'b0000000_100010000010;
      15'b011_100010010001 : VALUE=19'b0000000_100010000010;
      15'b011_100010010010 : VALUE=19'b0000000_100010000010;
      15'b011_100010010011 : VALUE=19'b0000000_100010000010;
      15'b011_100010010100 : VALUE=19'b0000000_100010000010;
      15'b011_100010010101 : VALUE=19'b0000000_100010000010;
      15'b011_100010010110 : VALUE=19'b0000000_100010000010;
      15'b011_100010010111 : VALUE=19'b0000000_100010000010;
      15'b011_100010011000 : VALUE=19'b0000000_100010000010;
      15'b011_100010011001 : VALUE=19'b0000000_100010000010;
      15'b011_100010011010 : VALUE=19'b0000000_100010000010;
      15'b011_100010011011 : VALUE=19'b0000000_100010000010;
      15'b011_100010011100 : VALUE=19'b0000000_100010000010;
      15'b011_100010011101 : VALUE=19'b0000000_100010000010;
      15'b011_100010011110 : VALUE=19'b0000000_100010000001;
      15'b011_100010011111 : VALUE=19'b0000000_100010000001;
      15'b011_100010100000 : VALUE=19'b0000000_100010000001;
      15'b011_100010100001 : VALUE=19'b0000000_100010000001;
      15'b011_100010100010 : VALUE=19'b0000000_100010000001;
      15'b011_100010100011 : VALUE=19'b0000000_100010000001;
      15'b011_100010100100 : VALUE=19'b0000000_100010000001;
      15'b011_100010100101 : VALUE=19'b0000000_100010000001;
      15'b011_100010100110 : VALUE=19'b0000000_100010000001;
      15'b011_100010100111 : VALUE=19'b0000000_100010000001;
      15'b011_100010101000 : VALUE=19'b0000000_100010000001;
      15'b011_100010101001 : VALUE=19'b0000000_100010000001;
      15'b011_100010101010 : VALUE=19'b0000000_100010000001;
      15'b011_100010101011 : VALUE=19'b0000000_100010000000;
      15'b011_100010101100 : VALUE=19'b0000000_100010000000;
      15'b011_100010101101 : VALUE=19'b0000000_100010000000;
      15'b011_100010101110 : VALUE=19'b0000000_100010000000;
      15'b011_100010101111 : VALUE=19'b0000000_100010000000;
      15'b011_100010110000 : VALUE=19'b0000000_100010000000;
      15'b011_100010110001 : VALUE=19'b0000000_100010000000;
      15'b011_100010110010 : VALUE=19'b0000000_100010000000;
      15'b011_100010110011 : VALUE=19'b0000000_100010000000;
      15'b011_100010110100 : VALUE=19'b0000000_100010000000;
      15'b011_100010110101 : VALUE=19'b0000000_100010000000;
      15'b011_100010110110 : VALUE=19'b0000000_100010000000;
      15'b011_100010110111 : VALUE=19'b0000000_100010000000;
      15'b011_100010111000 : VALUE=19'b0000000_100001111111;
      15'b011_100010111001 : VALUE=19'b0000000_100001111111;
      15'b011_100010111010 : VALUE=19'b0000000_100001111111;
      15'b011_100010111011 : VALUE=19'b0000000_100001111111;
      15'b011_100010111100 : VALUE=19'b0000000_100001111111;
      15'b011_100010111101 : VALUE=19'b0000000_100001111111;
      15'b011_100010111110 : VALUE=19'b0000000_100001111111;
      15'b011_100010111111 : VALUE=19'b0000000_100001111111;
      15'b011_100011000000 : VALUE=19'b0000000_100001111111;
      15'b011_100011000001 : VALUE=19'b0000000_100001111111;
      15'b011_100011000010 : VALUE=19'b0000000_100001111111;
      15'b011_100011000011 : VALUE=19'b0000000_100001111111;
      15'b011_100011000100 : VALUE=19'b0000000_100001111111;
      15'b011_100011000101 : VALUE=19'b0000000_100001111111;
      15'b011_100011000110 : VALUE=19'b0000000_100001111110;
      15'b011_100011000111 : VALUE=19'b0000000_100001111110;
      15'b011_100011001000 : VALUE=19'b0000000_100001111110;
      15'b011_100011001001 : VALUE=19'b0000000_100001111110;
      15'b011_100011001010 : VALUE=19'b0000000_100001111110;
      15'b011_100011001011 : VALUE=19'b0000000_100001111110;
      15'b011_100011001100 : VALUE=19'b0000000_100001111110;
      15'b011_100011001101 : VALUE=19'b0000000_100001111110;
      15'b011_100011001110 : VALUE=19'b0000000_100001111110;
      15'b011_100011001111 : VALUE=19'b0000000_100001111110;
      15'b011_100011010000 : VALUE=19'b0000000_100001111110;
      15'b011_100011010001 : VALUE=19'b0000000_100001111110;
      15'b011_100011010010 : VALUE=19'b0000000_100001111110;
      15'b011_100011010011 : VALUE=19'b0000000_100001111101;
      15'b011_100011010100 : VALUE=19'b0000000_100001111101;
      15'b011_100011010101 : VALUE=19'b0000000_100001111101;
      15'b011_100011010110 : VALUE=19'b0000000_100001111101;
      15'b011_100011010111 : VALUE=19'b0000000_100001111101;
      15'b011_100011011000 : VALUE=19'b0000000_100001111101;
      15'b011_100011011001 : VALUE=19'b0000000_100001111101;
      15'b011_100011011010 : VALUE=19'b0000000_100001111101;
      15'b011_100011011011 : VALUE=19'b0000000_100001111101;
      15'b011_100011011100 : VALUE=19'b0000000_100001111101;
      15'b011_100011011101 : VALUE=19'b0000000_100001111101;
      15'b011_100011011110 : VALUE=19'b0000000_100001111101;
      15'b011_100011011111 : VALUE=19'b0000000_100001111101;
      15'b011_100011100000 : VALUE=19'b0000000_100001111100;
      15'b011_100011100001 : VALUE=19'b0000000_100001111100;
      15'b011_100011100010 : VALUE=19'b0000000_100001111100;
      15'b011_100011100011 : VALUE=19'b0000000_100001111100;
      15'b011_100011100100 : VALUE=19'b0000000_100001111100;
      15'b011_100011100101 : VALUE=19'b0000000_100001111100;
      15'b011_100011100110 : VALUE=19'b0000000_100001111100;
      15'b011_100011100111 : VALUE=19'b0000000_100001111100;
      15'b011_100011101000 : VALUE=19'b0000000_100001111100;
      15'b011_100011101001 : VALUE=19'b0000000_100001111100;
      15'b011_100011101010 : VALUE=19'b0000000_100001111100;
      15'b011_100011101011 : VALUE=19'b0000000_100001111100;
      15'b011_100011101100 : VALUE=19'b0000000_100001111100;
      15'b011_100011101101 : VALUE=19'b0000000_100001111100;
      15'b011_100011101110 : VALUE=19'b0000000_100001111011;
      15'b011_100011101111 : VALUE=19'b0000000_100001111011;
      15'b011_100011110000 : VALUE=19'b0000000_100001111011;
      15'b011_100011110001 : VALUE=19'b0000000_100001111011;
      15'b011_100011110010 : VALUE=19'b0000000_100001111011;
      15'b011_100011110011 : VALUE=19'b0000000_100001111011;
      15'b011_100011110100 : VALUE=19'b0000000_100001111011;
      15'b011_100011110101 : VALUE=19'b0000000_100001111011;
      15'b011_100011110110 : VALUE=19'b0000000_100001111011;
      15'b011_100011110111 : VALUE=19'b0000000_100001111011;
      15'b011_100011111000 : VALUE=19'b0000000_100001111011;
      15'b011_100011111001 : VALUE=19'b0000000_100001111011;
      15'b011_100011111010 : VALUE=19'b0000000_100001111011;
      15'b011_100011111011 : VALUE=19'b0000000_100001111010;
      15'b011_100011111100 : VALUE=19'b0000000_100001111010;
      15'b011_100011111101 : VALUE=19'b0000000_100001111010;
      15'b011_100011111110 : VALUE=19'b0000000_100001111010;
      15'b011_100011111111 : VALUE=19'b0000000_100001111010;
      15'b011_100100000000 : VALUE=19'b0000000_100001111010;
      15'b011_100100000001 : VALUE=19'b0000000_100001111010;
      15'b011_100100000010 : VALUE=19'b0000000_100001111010;
      15'b011_100100000011 : VALUE=19'b0000000_100001111010;
      15'b011_100100000100 : VALUE=19'b0000000_100001111010;
      15'b011_100100000101 : VALUE=19'b0000000_100001111010;
      15'b011_100100000110 : VALUE=19'b0000000_100001111010;
      15'b011_100100000111 : VALUE=19'b0000000_100001111010;
      15'b011_100100001000 : VALUE=19'b0000000_100001111010;
      15'b011_100100001001 : VALUE=19'b0000000_100001111001;
      15'b011_100100001010 : VALUE=19'b0000000_100001111001;
      15'b011_100100001011 : VALUE=19'b0000000_100001111001;
      15'b011_100100001100 : VALUE=19'b0000000_100001111001;
      15'b011_100100001101 : VALUE=19'b0000000_100001111001;
      15'b011_100100001110 : VALUE=19'b0000000_100001111001;
      15'b011_100100001111 : VALUE=19'b0000000_100001111001;
      15'b011_100100010000 : VALUE=19'b0000000_100001111001;
      15'b011_100100010001 : VALUE=19'b0000000_100001111001;
      15'b011_100100010010 : VALUE=19'b0000000_100001111001;
      15'b011_100100010011 : VALUE=19'b0000000_100001111001;
      15'b011_100100010100 : VALUE=19'b0000000_100001111001;
      15'b011_100100010101 : VALUE=19'b0000000_100001111001;
      15'b011_100100010110 : VALUE=19'b0000000_100001111000;
      15'b011_100100010111 : VALUE=19'b0000000_100001111000;
      15'b011_100100011000 : VALUE=19'b0000000_100001111000;
      15'b011_100100011001 : VALUE=19'b0000000_100001111000;
      15'b011_100100011010 : VALUE=19'b0000000_100001111000;
      15'b011_100100011011 : VALUE=19'b0000000_100001111000;
      15'b011_100100011100 : VALUE=19'b0000000_100001111000;
      15'b011_100100011101 : VALUE=19'b0000000_100001111000;
      15'b011_100100011110 : VALUE=19'b0000000_100001111000;
      15'b011_100100011111 : VALUE=19'b0000000_100001111000;
      15'b011_100100100000 : VALUE=19'b0000000_100001111000;
      15'b011_100100100001 : VALUE=19'b0000000_100001111000;
      15'b011_100100100010 : VALUE=19'b0000000_100001111000;
      15'b011_100100100011 : VALUE=19'b0000000_100001111000;
      15'b011_100100100100 : VALUE=19'b0000000_100001110111;
      15'b011_100100100101 : VALUE=19'b0000000_100001110111;
      15'b011_100100100110 : VALUE=19'b0000000_100001110111;
      15'b011_100100100111 : VALUE=19'b0000000_100001110111;
      15'b011_100100101000 : VALUE=19'b0000000_100001110111;
      15'b011_100100101001 : VALUE=19'b0000000_100001110111;
      15'b011_100100101010 : VALUE=19'b0000000_100001110111;
      15'b011_100100101011 : VALUE=19'b0000000_100001110111;
      15'b011_100100101100 : VALUE=19'b0000000_100001110111;
      15'b011_100100101101 : VALUE=19'b0000000_100001110111;
      15'b011_100100101110 : VALUE=19'b0000000_100001110111;
      15'b011_100100101111 : VALUE=19'b0000000_100001110111;
      15'b011_100100110000 : VALUE=19'b0000000_100001110111;
      15'b011_100100110001 : VALUE=19'b0000000_100001110110;
      15'b011_100100110010 : VALUE=19'b0000000_100001110110;
      15'b011_100100110011 : VALUE=19'b0000000_100001110110;
      15'b011_100100110100 : VALUE=19'b0000000_100001110110;
      15'b011_100100110101 : VALUE=19'b0000000_100001110110;
      15'b011_100100110110 : VALUE=19'b0000000_100001110110;
      15'b011_100100110111 : VALUE=19'b0000000_100001110110;
      15'b011_100100111000 : VALUE=19'b0000000_100001110110;
      15'b011_100100111001 : VALUE=19'b0000000_100001110110;
      15'b011_100100111010 : VALUE=19'b0000000_100001110110;
      15'b011_100100111011 : VALUE=19'b0000000_100001110110;
      15'b011_100100111100 : VALUE=19'b0000000_100001110110;
      15'b011_100100111101 : VALUE=19'b0000000_100001110110;
      15'b011_100100111110 : VALUE=19'b0000000_100001110110;
      15'b011_100100111111 : VALUE=19'b0000000_100001110101;
      15'b011_100101000000 : VALUE=19'b0000000_100001110101;
      15'b011_100101000001 : VALUE=19'b0000000_100001110101;
      15'b011_100101000010 : VALUE=19'b0000000_100001110101;
      15'b011_100101000011 : VALUE=19'b0000000_100001110101;
      15'b011_100101000100 : VALUE=19'b0000000_100001110101;
      15'b011_100101000101 : VALUE=19'b0000000_100001110101;
      15'b011_100101000110 : VALUE=19'b0000000_100001110101;
      15'b011_100101000111 : VALUE=19'b0000000_100001110101;
      15'b011_100101001000 : VALUE=19'b0000000_100001110101;
      15'b011_100101001001 : VALUE=19'b0000000_100001110101;
      15'b011_100101001010 : VALUE=19'b0000000_100001110101;
      15'b011_100101001011 : VALUE=19'b0000000_100001110101;
      15'b011_100101001100 : VALUE=19'b0000000_100001110100;
      15'b011_100101001101 : VALUE=19'b0000000_100001110100;
      15'b011_100101001110 : VALUE=19'b0000000_100001110100;
      15'b011_100101001111 : VALUE=19'b0000000_100001110100;
      15'b011_100101010000 : VALUE=19'b0000000_100001110100;
      15'b011_100101010001 : VALUE=19'b0000000_100001110100;
      15'b011_100101010010 : VALUE=19'b0000000_100001110100;
      15'b011_100101010011 : VALUE=19'b0000000_100001110100;
      15'b011_100101010100 : VALUE=19'b0000000_100001110100;
      15'b011_100101010101 : VALUE=19'b0000000_100001110100;
      15'b011_100101010110 : VALUE=19'b0000000_100001110100;
      15'b011_100101010111 : VALUE=19'b0000000_100001110100;
      15'b011_100101011000 : VALUE=19'b0000000_100001110100;
      15'b011_100101011001 : VALUE=19'b0000000_100001110100;
      15'b011_100101011010 : VALUE=19'b0000000_100001110011;
      15'b011_100101011011 : VALUE=19'b0000000_100001110011;
      15'b011_100101011100 : VALUE=19'b0000000_100001110011;
      15'b011_100101011101 : VALUE=19'b0000000_100001110011;
      15'b011_100101011110 : VALUE=19'b0000000_100001110011;
      15'b011_100101011111 : VALUE=19'b0000000_100001110011;
      15'b011_100101100000 : VALUE=19'b0000000_100001110011;
      15'b011_100101100001 : VALUE=19'b0000000_100001110011;
      15'b011_100101100010 : VALUE=19'b0000000_100001110011;
      15'b011_100101100011 : VALUE=19'b0000000_100001110011;
      15'b011_100101100100 : VALUE=19'b0000000_100001110011;
      15'b011_100101100101 : VALUE=19'b0000000_100001110011;
      15'b011_100101100110 : VALUE=19'b0000000_100001110011;
      15'b011_100101100111 : VALUE=19'b0000000_100001110010;
      15'b011_100101101000 : VALUE=19'b0000000_100001110010;
      15'b011_100101101001 : VALUE=19'b0000000_100001110010;
      15'b011_100101101010 : VALUE=19'b0000000_100001110010;
      15'b011_100101101011 : VALUE=19'b0000000_100001110010;
      15'b011_100101101100 : VALUE=19'b0000000_100001110010;
      15'b011_100101101101 : VALUE=19'b0000000_100001110010;
      15'b011_100101101110 : VALUE=19'b0000000_100001110010;
      15'b011_100101101111 : VALUE=19'b0000000_100001110010;
      15'b011_100101110000 : VALUE=19'b0000000_100001110010;
      15'b011_100101110001 : VALUE=19'b0000000_100001110010;
      15'b011_100101110010 : VALUE=19'b0000000_100001110010;
      15'b011_100101110011 : VALUE=19'b0000000_100001110010;
      15'b011_100101110100 : VALUE=19'b0000000_100001110010;
      15'b011_100101110101 : VALUE=19'b0000000_100001110001;
      15'b011_100101110110 : VALUE=19'b0000000_100001110001;
      15'b011_100101110111 : VALUE=19'b0000000_100001110001;
      15'b011_100101111000 : VALUE=19'b0000000_100001110001;
      15'b011_100101111001 : VALUE=19'b0000000_100001110001;
      15'b011_100101111010 : VALUE=19'b0000000_100001110001;
      15'b011_100101111011 : VALUE=19'b0000000_100001110001;
      15'b011_100101111100 : VALUE=19'b0000000_100001110001;
      15'b011_100101111101 : VALUE=19'b0000000_100001110001;
      15'b011_100101111110 : VALUE=19'b0000000_100001110001;
      15'b011_100101111111 : VALUE=19'b0000000_100001110001;
      15'b011_100110000000 : VALUE=19'b0000000_100001110001;
      15'b011_100110000001 : VALUE=19'b0000000_100001110001;
      15'b011_100110000010 : VALUE=19'b0000000_100001110001;
      15'b011_100110000011 : VALUE=19'b0000000_100001110000;
      15'b011_100110000100 : VALUE=19'b0000000_100001110000;
      15'b011_100110000101 : VALUE=19'b0000000_100001110000;
      15'b011_100110000110 : VALUE=19'b0000000_100001110000;
      15'b011_100110000111 : VALUE=19'b0000000_100001110000;
      15'b011_100110001000 : VALUE=19'b0000000_100001110000;
      15'b011_100110001001 : VALUE=19'b0000000_100001110000;
      15'b011_100110001010 : VALUE=19'b0000000_100001110000;
      15'b011_100110001011 : VALUE=19'b0000000_100001110000;
      15'b011_100110001100 : VALUE=19'b0000000_100001110000;
      15'b011_100110001101 : VALUE=19'b0000000_100001110000;
      15'b011_100110001110 : VALUE=19'b0000000_100001110000;
      15'b011_100110001111 : VALUE=19'b0000000_100001110000;
      15'b011_100110010000 : VALUE=19'b0000000_100001101111;
      15'b011_100110010001 : VALUE=19'b0000000_100001101111;
      15'b011_100110010010 : VALUE=19'b0000000_100001101111;
      15'b011_100110010011 : VALUE=19'b0000000_100001101111;
      15'b011_100110010100 : VALUE=19'b0000000_100001101111;
      15'b011_100110010101 : VALUE=19'b0000000_100001101111;
      15'b011_100110010110 : VALUE=19'b0000000_100001101111;
      15'b011_100110010111 : VALUE=19'b0000000_100001101111;
      15'b011_100110011000 : VALUE=19'b0000000_100001101111;
      15'b011_100110011001 : VALUE=19'b0000000_100001101111;
      15'b011_100110011010 : VALUE=19'b0000000_100001101111;
      15'b011_100110011011 : VALUE=19'b0000000_100001101111;
      15'b011_100110011100 : VALUE=19'b0000000_100001101111;
      15'b011_100110011101 : VALUE=19'b0000000_100001101111;
      15'b011_100110011110 : VALUE=19'b0000000_100001101110;
      15'b011_100110011111 : VALUE=19'b0000000_100001101110;
      15'b011_100110100000 : VALUE=19'b0000000_100001101110;
      15'b011_100110100001 : VALUE=19'b0000000_100001101110;
      15'b011_100110100010 : VALUE=19'b0000000_100001101110;
      15'b011_100110100011 : VALUE=19'b0000000_100001101110;
      15'b011_100110100100 : VALUE=19'b0000000_100001101110;
      15'b011_100110100101 : VALUE=19'b0000000_100001101110;
      15'b011_100110100110 : VALUE=19'b0000000_100001101110;
      15'b011_100110100111 : VALUE=19'b0000000_100001101110;
      15'b011_100110101000 : VALUE=19'b0000000_100001101110;
      15'b011_100110101001 : VALUE=19'b0000000_100001101110;
      15'b011_100110101010 : VALUE=19'b0000000_100001101110;
      15'b011_100110101011 : VALUE=19'b0000000_100001101110;
      15'b011_100110101100 : VALUE=19'b0000000_100001101101;
      15'b011_100110101101 : VALUE=19'b0000000_100001101101;
      15'b011_100110101110 : VALUE=19'b0000000_100001101101;
      15'b011_100110101111 : VALUE=19'b0000000_100001101101;
      15'b011_100110110000 : VALUE=19'b0000000_100001101101;
      15'b011_100110110001 : VALUE=19'b0000000_100001101101;
      15'b011_100110110010 : VALUE=19'b0000000_100001101101;
      15'b011_100110110011 : VALUE=19'b0000000_100001101101;
      15'b011_100110110100 : VALUE=19'b0000000_100001101101;
      15'b011_100110110101 : VALUE=19'b0000000_100001101101;
      15'b011_100110110110 : VALUE=19'b0000000_100001101101;
      15'b011_100110110111 : VALUE=19'b0000000_100001101101;
      15'b011_100110111000 : VALUE=19'b0000000_100001101101;
      15'b011_100110111001 : VALUE=19'b0000000_100001101100;
      15'b011_100110111010 : VALUE=19'b0000000_100001101100;
      15'b011_100110111011 : VALUE=19'b0000000_100001101100;
      15'b011_100110111100 : VALUE=19'b0000000_100001101100;
      15'b011_100110111101 : VALUE=19'b0000000_100001101100;
      15'b011_100110111110 : VALUE=19'b0000000_100001101100;
      15'b011_100110111111 : VALUE=19'b0000000_100001101100;
      15'b011_100111000000 : VALUE=19'b0000000_100001101100;
      15'b011_100111000001 : VALUE=19'b0000000_100001101100;
      15'b011_100111000010 : VALUE=19'b0000000_100001101100;
      15'b011_100111000011 : VALUE=19'b0000000_100001101100;
      15'b011_100111000100 : VALUE=19'b0000000_100001101100;
      15'b011_100111000101 : VALUE=19'b0000000_100001101100;
      15'b011_100111000110 : VALUE=19'b0000000_100001101100;
      15'b011_100111000111 : VALUE=19'b0000000_100001101011;
      15'b011_100111001000 : VALUE=19'b0000000_100001101011;
      15'b011_100111001001 : VALUE=19'b0000000_100001101011;
      15'b011_100111001010 : VALUE=19'b0000000_100001101011;
      15'b011_100111001011 : VALUE=19'b0000000_100001101011;
      15'b011_100111001100 : VALUE=19'b0000000_100001101011;
      15'b011_100111001101 : VALUE=19'b0000000_100001101011;
      15'b011_100111001110 : VALUE=19'b0000000_100001101011;
      15'b011_100111001111 : VALUE=19'b0000000_100001101011;
      15'b011_100111010000 : VALUE=19'b0000000_100001101011;
      15'b011_100111010001 : VALUE=19'b0000000_100001101011;
      15'b011_100111010010 : VALUE=19'b0000000_100001101011;
      15'b011_100111010011 : VALUE=19'b0000000_100001101011;
      15'b011_100111010100 : VALUE=19'b0000000_100001101011;
      15'b011_100111010101 : VALUE=19'b0000000_100001101010;
      15'b011_100111010110 : VALUE=19'b0000000_100001101010;
      15'b011_100111010111 : VALUE=19'b0000000_100001101010;
      15'b011_100111011000 : VALUE=19'b0000000_100001101010;
      15'b011_100111011001 : VALUE=19'b0000000_100001101010;
      15'b011_100111011010 : VALUE=19'b0000000_100001101010;
      15'b011_100111011011 : VALUE=19'b0000000_100001101010;
      15'b011_100111011100 : VALUE=19'b0000000_100001101010;
      15'b011_100111011101 : VALUE=19'b0000000_100001101010;
      15'b011_100111011110 : VALUE=19'b0000000_100001101010;
      15'b011_100111011111 : VALUE=19'b0000000_100001101010;
      15'b011_100111100000 : VALUE=19'b0000000_100001101010;
      15'b011_100111100001 : VALUE=19'b0000000_100001101010;
      15'b011_100111100010 : VALUE=19'b0000000_100001101010;
      15'b011_100111100011 : VALUE=19'b0000000_100001101001;
      15'b011_100111100100 : VALUE=19'b0000000_100001101001;
      15'b011_100111100101 : VALUE=19'b0000000_100001101001;
      15'b011_100111100110 : VALUE=19'b0000000_100001101001;
      15'b011_100111100111 : VALUE=19'b0000000_100001101001;
      15'b011_100111101000 : VALUE=19'b0000000_100001101001;
      15'b011_100111101001 : VALUE=19'b0000000_100001101001;
      15'b011_100111101010 : VALUE=19'b0000000_100001101001;
      15'b011_100111101011 : VALUE=19'b0000000_100001101001;
      15'b011_100111101100 : VALUE=19'b0000000_100001101001;
      15'b011_100111101101 : VALUE=19'b0000000_100001101001;
      15'b011_100111101110 : VALUE=19'b0000000_100001101001;
      15'b011_100111101111 : VALUE=19'b0000000_100001101001;
      15'b011_100111110000 : VALUE=19'b0000000_100001101000;
      15'b011_100111110001 : VALUE=19'b0000000_100001101000;
      15'b011_100111110010 : VALUE=19'b0000000_100001101000;
      15'b011_100111110011 : VALUE=19'b0000000_100001101000;
      15'b011_100111110100 : VALUE=19'b0000000_100001101000;
      15'b011_100111110101 : VALUE=19'b0000000_100001101000;
      15'b011_100111110110 : VALUE=19'b0000000_100001101000;
      15'b011_100111110111 : VALUE=19'b0000000_100001101000;
      15'b011_100111111000 : VALUE=19'b0000000_100001101000;
      15'b011_100111111001 : VALUE=19'b0000000_100001101000;
      15'b011_100111111010 : VALUE=19'b0000000_100001101000;
      15'b011_100111111011 : VALUE=19'b0000000_100001101000;
      15'b011_100111111100 : VALUE=19'b0000000_100001101000;
      15'b011_100111111101 : VALUE=19'b0000000_100001101000;
      15'b011_100111111110 : VALUE=19'b0000000_100001100111;
      15'b011_100111111111 : VALUE=19'b0000000_100001100111;
      15'b011_101000000000 : VALUE=19'b0000000_100001100111;
      15'b011_101000000001 : VALUE=19'b0000000_100001100111;
      15'b011_101000000010 : VALUE=19'b0000000_100001100111;
      15'b011_101000000011 : VALUE=19'b0000000_100001100111;
      15'b011_101000000100 : VALUE=19'b0000000_100001100111;
      15'b011_101000000101 : VALUE=19'b0000000_100001100111;
      15'b011_101000000110 : VALUE=19'b0000000_100001100111;
      15'b011_101000000111 : VALUE=19'b0000000_100001100111;
      15'b011_101000001000 : VALUE=19'b0000000_100001100111;
      15'b011_101000001001 : VALUE=19'b0000000_100001100111;
      15'b011_101000001010 : VALUE=19'b0000000_100001100111;
      15'b011_101000001011 : VALUE=19'b0000000_100001100111;
      15'b011_101000001100 : VALUE=19'b0000000_100001100110;
      15'b011_101000001101 : VALUE=19'b0000000_100001100110;
      15'b011_101000001110 : VALUE=19'b0000000_100001100110;
      15'b011_101000001111 : VALUE=19'b0000000_100001100110;
      15'b011_101000010000 : VALUE=19'b0000000_100001100110;
      15'b011_101000010001 : VALUE=19'b0000000_100001100110;
      15'b011_101000010010 : VALUE=19'b0000000_100001100110;
      15'b011_101000010011 : VALUE=19'b0000000_100001100110;
      15'b011_101000010100 : VALUE=19'b0000000_100001100110;
      15'b011_101000010101 : VALUE=19'b0000000_100001100110;
      15'b011_101000010110 : VALUE=19'b0000000_100001100110;
      15'b011_101000010111 : VALUE=19'b0000000_100001100110;
      15'b011_101000011000 : VALUE=19'b0000000_100001100110;
      15'b011_101000011001 : VALUE=19'b0000000_100001100110;
      15'b011_101000011010 : VALUE=19'b0000000_100001100101;
      15'b011_101000011011 : VALUE=19'b0000000_100001100101;
      15'b011_101000011100 : VALUE=19'b0000000_100001100101;
      15'b011_101000011101 : VALUE=19'b0000000_100001100101;
      15'b011_101000011110 : VALUE=19'b0000000_100001100101;
      15'b011_101000011111 : VALUE=19'b0000000_100001100101;
      15'b011_101000100000 : VALUE=19'b0000000_100001100101;
      15'b011_101000100001 : VALUE=19'b0000000_100001100101;
      15'b011_101000100010 : VALUE=19'b0000000_100001100101;
      15'b011_101000100011 : VALUE=19'b0000000_100001100101;
      15'b011_101000100100 : VALUE=19'b0000000_100001100101;
      15'b011_101000100101 : VALUE=19'b0000000_100001100101;
      15'b011_101000100110 : VALUE=19'b0000000_100001100101;
      15'b011_101000100111 : VALUE=19'b0000000_100001100101;
      15'b011_101000101000 : VALUE=19'b0000000_100001100100;
      15'b011_101000101001 : VALUE=19'b0000000_100001100100;
      15'b011_101000101010 : VALUE=19'b0000000_100001100100;
      15'b011_101000101011 : VALUE=19'b0000000_100001100100;
      15'b011_101000101100 : VALUE=19'b0000000_100001100100;
      15'b011_101000101101 : VALUE=19'b0000000_100001100100;
      15'b011_101000101110 : VALUE=19'b0000000_100001100100;
      15'b011_101000101111 : VALUE=19'b0000000_100001100100;
      15'b011_101000110000 : VALUE=19'b0000000_100001100100;
      15'b011_101000110001 : VALUE=19'b0000000_100001100100;
      15'b011_101000110010 : VALUE=19'b0000000_100001100100;
      15'b011_101000110011 : VALUE=19'b0000000_100001100100;
      15'b011_101000110100 : VALUE=19'b0000000_100001100100;
      15'b011_101000110101 : VALUE=19'b0000000_100001100011;
      15'b011_101000110110 : VALUE=19'b0000000_100001100011;
      15'b011_101000110111 : VALUE=19'b0000000_100001100011;
      15'b011_101000111000 : VALUE=19'b0000000_100001100011;
      15'b011_101000111001 : VALUE=19'b0000000_100001100011;
      15'b011_101000111010 : VALUE=19'b0000000_100001100011;
      15'b011_101000111011 : VALUE=19'b0000000_100001100011;
      15'b011_101000111100 : VALUE=19'b0000000_100001100011;
      15'b011_101000111101 : VALUE=19'b0000000_100001100011;
      15'b011_101000111110 : VALUE=19'b0000000_100001100011;
      15'b011_101000111111 : VALUE=19'b0000000_100001100011;
      15'b011_101001000000 : VALUE=19'b0000000_100001100011;
      15'b011_101001000001 : VALUE=19'b0000000_100001100011;
      15'b011_101001000010 : VALUE=19'b0000000_100001100011;
      15'b011_101001000011 : VALUE=19'b0000000_100001100010;
      15'b011_101001000100 : VALUE=19'b0000000_100001100010;
      15'b011_101001000101 : VALUE=19'b0000000_100001100010;
      15'b011_101001000110 : VALUE=19'b0000000_100001100010;
      15'b011_101001000111 : VALUE=19'b0000000_100001100010;
      15'b011_101001001000 : VALUE=19'b0000000_100001100010;
      15'b011_101001001001 : VALUE=19'b0000000_100001100010;
      15'b011_101001001010 : VALUE=19'b0000000_100001100010;
      15'b011_101001001011 : VALUE=19'b0000000_100001100010;
      15'b011_101001001100 : VALUE=19'b0000000_100001100010;
      15'b011_101001001101 : VALUE=19'b0000000_100001100010;
      15'b011_101001001110 : VALUE=19'b0000000_100001100010;
      15'b011_101001001111 : VALUE=19'b0000000_100001100010;
      15'b011_101001010000 : VALUE=19'b0000000_100001100010;
      15'b011_101001010001 : VALUE=19'b0000000_100001100001;
      15'b011_101001010010 : VALUE=19'b0000000_100001100001;
      15'b011_101001010011 : VALUE=19'b0000000_100001100001;
      15'b011_101001010100 : VALUE=19'b0000000_100001100001;
      15'b011_101001010101 : VALUE=19'b0000000_100001100001;
      15'b011_101001010110 : VALUE=19'b0000000_100001100001;
      15'b011_101001010111 : VALUE=19'b0000000_100001100001;
      15'b011_101001011000 : VALUE=19'b0000000_100001100001;
      15'b011_101001011001 : VALUE=19'b0000000_100001100001;
      15'b011_101001011010 : VALUE=19'b0000000_100001100001;
      15'b011_101001011011 : VALUE=19'b0000000_100001100001;
      15'b011_101001011100 : VALUE=19'b0000000_100001100001;
      15'b011_101001011101 : VALUE=19'b0000000_100001100001;
      15'b011_101001011110 : VALUE=19'b0000000_100001100001;
      15'b011_101001011111 : VALUE=19'b0000000_100001100000;
      15'b011_101001100000 : VALUE=19'b0000000_100001100000;
      15'b011_101001100001 : VALUE=19'b0000000_100001100000;
      15'b011_101001100010 : VALUE=19'b0000000_100001100000;
      15'b011_101001100011 : VALUE=19'b0000000_100001100000;
      15'b011_101001100100 : VALUE=19'b0000000_100001100000;
      15'b011_101001100101 : VALUE=19'b0000000_100001100000;
      15'b011_101001100110 : VALUE=19'b0000000_100001100000;
      15'b011_101001100111 : VALUE=19'b0000000_100001100000;
      15'b011_101001101000 : VALUE=19'b0000000_100001100000;
      15'b011_101001101001 : VALUE=19'b0000000_100001100000;
      15'b011_101001101010 : VALUE=19'b0000000_100001100000;
      15'b011_101001101011 : VALUE=19'b0000000_100001100000;
      15'b011_101001101100 : VALUE=19'b0000000_100001100000;
      15'b011_101001101101 : VALUE=19'b0000000_100001011111;
      15'b011_101001101110 : VALUE=19'b0000000_100001011111;
      15'b011_101001101111 : VALUE=19'b0000000_100001011111;
      15'b011_101001110000 : VALUE=19'b0000000_100001011111;
      15'b011_101001110001 : VALUE=19'b0000000_100001011111;
      15'b011_101001110010 : VALUE=19'b0000000_100001011111;
      15'b011_101001110011 : VALUE=19'b0000000_100001011111;
      15'b011_101001110100 : VALUE=19'b0000000_100001011111;
      15'b011_101001110101 : VALUE=19'b0000000_100001011111;
      15'b011_101001110110 : VALUE=19'b0000000_100001011111;
      15'b011_101001110111 : VALUE=19'b0000000_100001011111;
      15'b011_101001111000 : VALUE=19'b0000000_100001011111;
      15'b011_101001111001 : VALUE=19'b0000000_100001011111;
      15'b011_101001111010 : VALUE=19'b0000000_100001011111;
      15'b011_101001111011 : VALUE=19'b0000000_100001011110;
      15'b011_101001111100 : VALUE=19'b0000000_100001011110;
      15'b011_101001111101 : VALUE=19'b0000000_100001011110;
      15'b011_101001111110 : VALUE=19'b0000000_100001011110;
      15'b011_101001111111 : VALUE=19'b0000000_100001011110;
      15'b011_101010000000 : VALUE=19'b0000000_100001011110;
      15'b011_101010000001 : VALUE=19'b0000000_100001011110;
      15'b011_101010000010 : VALUE=19'b0000000_100001011110;
      15'b011_101010000011 : VALUE=19'b0000000_100001011110;
      15'b011_101010000100 : VALUE=19'b0000000_100001011110;
      15'b011_101010000101 : VALUE=19'b0000000_100001011110;
      15'b011_101010000110 : VALUE=19'b0000000_100001011110;
      15'b011_101010000111 : VALUE=19'b0000000_100001011110;
      15'b011_101010001000 : VALUE=19'b0000000_100001011110;
      15'b011_101010001001 : VALUE=19'b0000000_100001011101;
      15'b011_101010001010 : VALUE=19'b0000000_100001011101;
      15'b011_101010001011 : VALUE=19'b0000000_100001011101;
      15'b011_101010001100 : VALUE=19'b0000000_100001011101;
      15'b011_101010001101 : VALUE=19'b0000000_100001011101;
      15'b011_101010001110 : VALUE=19'b0000000_100001011101;
      15'b011_101010001111 : VALUE=19'b0000000_100001011101;
      15'b011_101010010000 : VALUE=19'b0000000_100001011101;
      15'b011_101010010001 : VALUE=19'b0000000_100001011101;
      15'b011_101010010010 : VALUE=19'b0000000_100001011101;
      15'b011_101010010011 : VALUE=19'b0000000_100001011101;
      15'b011_101010010100 : VALUE=19'b0000000_100001011101;
      15'b011_101010010101 : VALUE=19'b0000000_100001011101;
      15'b011_101010010110 : VALUE=19'b0000000_100001011101;
      15'b011_101010010111 : VALUE=19'b0000000_100001011100;
      15'b011_101010011000 : VALUE=19'b0000000_100001011100;
      15'b011_101010011001 : VALUE=19'b0000000_100001011100;
      15'b011_101010011010 : VALUE=19'b0000000_100001011100;
      15'b011_101010011011 : VALUE=19'b0000000_100001011100;
      15'b011_101010011100 : VALUE=19'b0000000_100001011100;
      15'b011_101010011101 : VALUE=19'b0000000_100001011100;
      15'b011_101010011110 : VALUE=19'b0000000_100001011100;
      15'b011_101010011111 : VALUE=19'b0000000_100001011100;
      15'b011_101010100000 : VALUE=19'b0000000_100001011100;
      15'b011_101010100001 : VALUE=19'b0000000_100001011100;
      15'b011_101010100010 : VALUE=19'b0000000_100001011100;
      15'b011_101010100011 : VALUE=19'b0000000_100001011100;
      15'b011_101010100100 : VALUE=19'b0000000_100001011100;
      15'b011_101010100101 : VALUE=19'b0000000_100001011011;
      15'b011_101010100110 : VALUE=19'b0000000_100001011011;
      15'b011_101010100111 : VALUE=19'b0000000_100001011011;
      15'b011_101010101000 : VALUE=19'b0000000_100001011011;
      15'b011_101010101001 : VALUE=19'b0000000_100001011011;
      15'b011_101010101010 : VALUE=19'b0000000_100001011011;
      15'b011_101010101011 : VALUE=19'b0000000_100001011011;
      15'b011_101010101100 : VALUE=19'b0000000_100001011011;
      15'b011_101010101101 : VALUE=19'b0000000_100001011011;
      15'b011_101010101110 : VALUE=19'b0000000_100001011011;
      15'b011_101010101111 : VALUE=19'b0000000_100001011011;
      15'b011_101010110000 : VALUE=19'b0000000_100001011011;
      15'b011_101010110001 : VALUE=19'b0000000_100001011011;
      15'b011_101010110010 : VALUE=19'b0000000_100001011011;
      15'b011_101010110011 : VALUE=19'b0000000_100001011010;
      15'b011_101010110100 : VALUE=19'b0000000_100001011010;
      15'b011_101010110101 : VALUE=19'b0000000_100001011010;
      15'b011_101010110110 : VALUE=19'b0000000_100001011010;
      15'b011_101010110111 : VALUE=19'b0000000_100001011010;
      15'b011_101010111000 : VALUE=19'b0000000_100001011010;
      15'b011_101010111001 : VALUE=19'b0000000_100001011010;
      15'b011_101010111010 : VALUE=19'b0000000_100001011010;
      15'b011_101010111011 : VALUE=19'b0000000_100001011010;
      15'b011_101010111100 : VALUE=19'b0000000_100001011010;
      15'b011_101010111101 : VALUE=19'b0000000_100001011010;
      15'b011_101010111110 : VALUE=19'b0000000_100001011010;
      15'b011_101010111111 : VALUE=19'b0000000_100001011010;
      15'b011_101011000000 : VALUE=19'b0000000_100001011010;
      15'b011_101011000001 : VALUE=19'b0000000_100001011001;
      15'b011_101011000010 : VALUE=19'b0000000_100001011001;
      15'b011_101011000011 : VALUE=19'b0000000_100001011001;
      15'b011_101011000100 : VALUE=19'b0000000_100001011001;
      15'b011_101011000101 : VALUE=19'b0000000_100001011001;
      15'b011_101011000110 : VALUE=19'b0000000_100001011001;
      15'b011_101011000111 : VALUE=19'b0000000_100001011001;
      15'b011_101011001000 : VALUE=19'b0000000_100001011001;
      15'b011_101011001001 : VALUE=19'b0000000_100001011001;
      15'b011_101011001010 : VALUE=19'b0000000_100001011001;
      15'b011_101011001011 : VALUE=19'b0000000_100001011001;
      15'b011_101011001100 : VALUE=19'b0000000_100001011001;
      15'b011_101011001101 : VALUE=19'b0000000_100001011001;
      15'b011_101011001110 : VALUE=19'b0000000_100001011001;
      15'b011_101011001111 : VALUE=19'b0000000_100001011000;
      15'b011_101011010000 : VALUE=19'b0000000_100001011000;
      15'b011_101011010001 : VALUE=19'b0000000_100001011000;
      15'b011_101011010010 : VALUE=19'b0000000_100001011000;
      15'b011_101011010011 : VALUE=19'b0000000_100001011000;
      15'b011_101011010100 : VALUE=19'b0000000_100001011000;
      15'b011_101011010101 : VALUE=19'b0000000_100001011000;
      15'b011_101011010110 : VALUE=19'b0000000_100001011000;
      15'b011_101011010111 : VALUE=19'b0000000_100001011000;
      15'b011_101011011000 : VALUE=19'b0000000_100001011000;
      15'b011_101011011001 : VALUE=19'b0000000_100001011000;
      15'b011_101011011010 : VALUE=19'b0000000_100001011000;
      15'b011_101011011011 : VALUE=19'b0000000_100001011000;
      15'b011_101011011100 : VALUE=19'b0000000_100001011000;
      15'b011_101011011101 : VALUE=19'b0000000_100001010111;
      15'b011_101011011110 : VALUE=19'b0000000_100001010111;
      15'b011_101011011111 : VALUE=19'b0000000_100001010111;
      15'b011_101011100000 : VALUE=19'b0000000_100001010111;
      15'b011_101011100001 : VALUE=19'b0000000_100001010111;
      15'b011_101011100010 : VALUE=19'b0000000_100001010111;
      15'b011_101011100011 : VALUE=19'b0000000_100001010111;
      15'b011_101011100100 : VALUE=19'b0000000_100001010111;
      15'b011_101011100101 : VALUE=19'b0000000_100001010111;
      15'b011_101011100110 : VALUE=19'b0000000_100001010111;
      15'b011_101011100111 : VALUE=19'b0000000_100001010111;
      15'b011_101011101000 : VALUE=19'b0000000_100001010111;
      15'b011_101011101001 : VALUE=19'b0000000_100001010111;
      15'b011_101011101010 : VALUE=19'b0000000_100001010111;
      15'b011_101011101011 : VALUE=19'b0000000_100001010110;
      15'b011_101011101100 : VALUE=19'b0000000_100001010110;
      15'b011_101011101101 : VALUE=19'b0000000_100001010110;
      15'b011_101011101110 : VALUE=19'b0000000_100001010110;
      15'b011_101011101111 : VALUE=19'b0000000_100001010110;
      15'b011_101011110000 : VALUE=19'b0000000_100001010110;
      15'b011_101011110001 : VALUE=19'b0000000_100001010110;
      15'b011_101011110010 : VALUE=19'b0000000_100001010110;
      15'b011_101011110011 : VALUE=19'b0000000_100001010110;
      15'b011_101011110100 : VALUE=19'b0000000_100001010110;
      15'b011_101011110101 : VALUE=19'b0000000_100001010110;
      15'b011_101011110110 : VALUE=19'b0000000_100001010110;
      15'b011_101011110111 : VALUE=19'b0000000_100001010110;
      15'b011_101011111000 : VALUE=19'b0000000_100001010110;
      15'b011_101011111001 : VALUE=19'b0000000_100001010110;
      15'b011_101011111010 : VALUE=19'b0000000_100001010101;
      15'b011_101011111011 : VALUE=19'b0000000_100001010101;
      15'b011_101011111100 : VALUE=19'b0000000_100001010101;
      15'b011_101011111101 : VALUE=19'b0000000_100001010101;
      15'b011_101011111110 : VALUE=19'b0000000_100001010101;
      15'b011_101011111111 : VALUE=19'b0000000_100001010101;
      15'b011_101100000000 : VALUE=19'b0000000_100001010101;
      15'b011_101100000001 : VALUE=19'b0000000_100001010101;
      15'b011_101100000010 : VALUE=19'b0000000_100001010101;
      15'b011_101100000011 : VALUE=19'b0000000_100001010101;
      15'b011_101100000100 : VALUE=19'b0000000_100001010101;
      15'b011_101100000101 : VALUE=19'b0000000_100001010101;
      15'b011_101100000110 : VALUE=19'b0000000_100001010101;
      15'b011_101100000111 : VALUE=19'b0000000_100001010101;
      15'b011_101100001000 : VALUE=19'b0000000_100001010100;
      15'b011_101100001001 : VALUE=19'b0000000_100001010100;
      15'b011_101100001010 : VALUE=19'b0000000_100001010100;
      15'b011_101100001011 : VALUE=19'b0000000_100001010100;
      15'b011_101100001100 : VALUE=19'b0000000_100001010100;
      15'b011_101100001101 : VALUE=19'b0000000_100001010100;
      15'b011_101100001110 : VALUE=19'b0000000_100001010100;
      15'b011_101100001111 : VALUE=19'b0000000_100001010100;
      15'b011_101100010000 : VALUE=19'b0000000_100001010100;
      15'b011_101100010001 : VALUE=19'b0000000_100001010100;
      15'b011_101100010010 : VALUE=19'b0000000_100001010100;
      15'b011_101100010011 : VALUE=19'b0000000_100001010100;
      15'b011_101100010100 : VALUE=19'b0000000_100001010100;
      15'b011_101100010101 : VALUE=19'b0000000_100001010100;
      15'b011_101100010110 : VALUE=19'b0000000_100001010011;
      15'b011_101100010111 : VALUE=19'b0000000_100001010011;
      15'b011_101100011000 : VALUE=19'b0000000_100001010011;
      15'b011_101100011001 : VALUE=19'b0000000_100001010011;
      15'b011_101100011010 : VALUE=19'b0000000_100001010011;
      15'b011_101100011011 : VALUE=19'b0000000_100001010011;
      15'b011_101100011100 : VALUE=19'b0000000_100001010011;
      15'b011_101100011101 : VALUE=19'b0000000_100001010011;
      15'b011_101100011110 : VALUE=19'b0000000_100001010011;
      15'b011_101100011111 : VALUE=19'b0000000_100001010011;
      15'b011_101100100000 : VALUE=19'b0000000_100001010011;
      15'b011_101100100001 : VALUE=19'b0000000_100001010011;
      15'b011_101100100010 : VALUE=19'b0000000_100001010011;
      15'b011_101100100011 : VALUE=19'b0000000_100001010011;
      15'b011_101100100100 : VALUE=19'b0000000_100001010010;
      15'b011_101100100101 : VALUE=19'b0000000_100001010010;
      15'b011_101100100110 : VALUE=19'b0000000_100001010010;
      15'b011_101100100111 : VALUE=19'b0000000_100001010010;
      15'b011_101100101000 : VALUE=19'b0000000_100001010010;
      15'b011_101100101001 : VALUE=19'b0000000_100001010010;
      15'b011_101100101010 : VALUE=19'b0000000_100001010010;
      15'b011_101100101011 : VALUE=19'b0000000_100001010010;
      15'b011_101100101100 : VALUE=19'b0000000_100001010010;
      15'b011_101100101101 : VALUE=19'b0000000_100001010010;
      15'b011_101100101110 : VALUE=19'b0000000_100001010010;
      15'b011_101100101111 : VALUE=19'b0000000_100001010010;
      15'b011_101100110000 : VALUE=19'b0000000_100001010010;
      15'b011_101100110001 : VALUE=19'b0000000_100001010010;
      15'b011_101100110010 : VALUE=19'b0000000_100001010001;
      15'b011_101100110011 : VALUE=19'b0000000_100001010001;
      15'b011_101100110100 : VALUE=19'b0000000_100001010001;
      15'b011_101100110101 : VALUE=19'b0000000_100001010001;
      15'b011_101100110110 : VALUE=19'b0000000_100001010001;
      15'b011_101100110111 : VALUE=19'b0000000_100001010001;
      15'b011_101100111000 : VALUE=19'b0000000_100001010001;
      15'b011_101100111001 : VALUE=19'b0000000_100001010001;
      15'b011_101100111010 : VALUE=19'b0000000_100001010001;
      15'b011_101100111011 : VALUE=19'b0000000_100001010001;
      15'b011_101100111100 : VALUE=19'b0000000_100001010001;
      15'b011_101100111101 : VALUE=19'b0000000_100001010001;
      15'b011_101100111110 : VALUE=19'b0000000_100001010001;
      15'b011_101100111111 : VALUE=19'b0000000_100001010001;
      15'b011_101101000000 : VALUE=19'b0000000_100001010001;
      15'b011_101101000001 : VALUE=19'b0000000_100001010000;
      15'b011_101101000010 : VALUE=19'b0000000_100001010000;
      15'b011_101101000011 : VALUE=19'b0000000_100001010000;
      15'b011_101101000100 : VALUE=19'b0000000_100001010000;
      15'b011_101101000101 : VALUE=19'b0000000_100001010000;
      15'b011_101101000110 : VALUE=19'b0000000_100001010000;
      15'b011_101101000111 : VALUE=19'b0000000_100001010000;
      15'b011_101101001000 : VALUE=19'b0000000_100001010000;
      15'b011_101101001001 : VALUE=19'b0000000_100001010000;
      15'b011_101101001010 : VALUE=19'b0000000_100001010000;
      15'b011_101101001011 : VALUE=19'b0000000_100001010000;
      15'b011_101101001100 : VALUE=19'b0000000_100001010000;
      15'b011_101101001101 : VALUE=19'b0000000_100001010000;
      15'b011_101101001110 : VALUE=19'b0000000_100001010000;
      15'b011_101101001111 : VALUE=19'b0000000_100001001111;
      15'b011_101101010000 : VALUE=19'b0000000_100001001111;
      15'b011_101101010001 : VALUE=19'b0000000_100001001111;
      15'b011_101101010010 : VALUE=19'b0000000_100001001111;
      15'b011_101101010011 : VALUE=19'b0000000_100001001111;
      15'b011_101101010100 : VALUE=19'b0000000_100001001111;
      15'b011_101101010101 : VALUE=19'b0000000_100001001111;
      15'b011_101101010110 : VALUE=19'b0000000_100001001111;
      15'b011_101101010111 : VALUE=19'b0000000_100001001111;
      15'b011_101101011000 : VALUE=19'b0000000_100001001111;
      15'b011_101101011001 : VALUE=19'b0000000_100001001111;
      15'b011_101101011010 : VALUE=19'b0000000_100001001111;
      15'b011_101101011011 : VALUE=19'b0000000_100001001111;
      15'b011_101101011100 : VALUE=19'b0000000_100001001111;
      15'b011_101101011101 : VALUE=19'b0000000_100001001110;
      15'b011_101101011110 : VALUE=19'b0000000_100001001110;
      15'b011_101101011111 : VALUE=19'b0000000_100001001110;
      15'b011_101101100000 : VALUE=19'b0000000_100001001110;
      15'b011_101101100001 : VALUE=19'b0000000_100001001110;
      15'b011_101101100010 : VALUE=19'b0000000_100001001110;
      15'b011_101101100011 : VALUE=19'b0000000_100001001110;
      15'b011_101101100100 : VALUE=19'b0000000_100001001110;
      15'b011_101101100101 : VALUE=19'b0000000_100001001110;
      15'b011_101101100110 : VALUE=19'b0000000_100001001110;
      15'b011_101101100111 : VALUE=19'b0000000_100001001110;
      15'b011_101101101000 : VALUE=19'b0000000_100001001110;
      15'b011_101101101001 : VALUE=19'b0000000_100001001110;
      15'b011_101101101010 : VALUE=19'b0000000_100001001110;
      15'b011_101101101011 : VALUE=19'b0000000_100001001101;
      15'b011_101101101100 : VALUE=19'b0000000_100001001101;
      15'b011_101101101101 : VALUE=19'b0000000_100001001101;
      15'b011_101101101110 : VALUE=19'b0000000_100001001101;
      15'b011_101101101111 : VALUE=19'b0000000_100001001101;
      15'b011_101101110000 : VALUE=19'b0000000_100001001101;
      15'b011_101101110001 : VALUE=19'b0000000_100001001101;
      15'b011_101101110010 : VALUE=19'b0000000_100001001101;
      15'b011_101101110011 : VALUE=19'b0000000_100001001101;
      15'b011_101101110100 : VALUE=19'b0000000_100001001101;
      15'b011_101101110101 : VALUE=19'b0000000_100001001101;
      15'b011_101101110110 : VALUE=19'b0000000_100001001101;
      15'b011_101101110111 : VALUE=19'b0000000_100001001101;
      15'b011_101101111000 : VALUE=19'b0000000_100001001101;
      15'b011_101101111001 : VALUE=19'b0000000_100001001101;
      15'b011_101101111010 : VALUE=19'b0000000_100001001100;
      15'b011_101101111011 : VALUE=19'b0000000_100001001100;
      15'b011_101101111100 : VALUE=19'b0000000_100001001100;
      15'b011_101101111101 : VALUE=19'b0000000_100001001100;
      15'b011_101101111110 : VALUE=19'b0000000_100001001100;
      15'b011_101101111111 : VALUE=19'b0000000_100001001100;
      15'b011_101110000000 : VALUE=19'b0000000_100001001100;
      15'b011_101110000001 : VALUE=19'b0000000_100001001100;
      15'b011_101110000010 : VALUE=19'b0000000_100001001100;
      15'b011_101110000011 : VALUE=19'b0000000_100001001100;
      15'b011_101110000100 : VALUE=19'b0000000_100001001100;
      15'b011_101110000101 : VALUE=19'b0000000_100001001100;
      15'b011_101110000110 : VALUE=19'b0000000_100001001100;
      15'b011_101110000111 : VALUE=19'b0000000_100001001100;
      15'b011_101110001000 : VALUE=19'b0000000_100001001011;
      15'b011_101110001001 : VALUE=19'b0000000_100001001011;
      15'b011_101110001010 : VALUE=19'b0000000_100001001011;
      15'b011_101110001011 : VALUE=19'b0000000_100001001011;
      15'b011_101110001100 : VALUE=19'b0000000_100001001011;
      15'b011_101110001101 : VALUE=19'b0000000_100001001011;
      15'b011_101110001110 : VALUE=19'b0000000_100001001011;
      15'b011_101110001111 : VALUE=19'b0000000_100001001011;
      15'b011_101110010000 : VALUE=19'b0000000_100001001011;
      15'b011_101110010001 : VALUE=19'b0000000_100001001011;
      15'b011_101110010010 : VALUE=19'b0000000_100001001011;
      15'b011_101110010011 : VALUE=19'b0000000_100001001011;
      15'b011_101110010100 : VALUE=19'b0000000_100001001011;
      15'b011_101110010101 : VALUE=19'b0000000_100001001011;
      15'b011_101110010110 : VALUE=19'b0000000_100001001011;
      15'b011_101110010111 : VALUE=19'b0000000_100001001010;
      15'b011_101110011000 : VALUE=19'b0000000_100001001010;
      15'b011_101110011001 : VALUE=19'b0000000_100001001010;
      15'b011_101110011010 : VALUE=19'b0000000_100001001010;
      15'b011_101110011011 : VALUE=19'b0000000_100001001010;
      15'b011_101110011100 : VALUE=19'b0000000_100001001010;
      15'b011_101110011101 : VALUE=19'b0000000_100001001010;
      15'b011_101110011110 : VALUE=19'b0000000_100001001010;
      15'b011_101110011111 : VALUE=19'b0000000_100001001010;
      15'b011_101110100000 : VALUE=19'b0000000_100001001010;
      15'b011_101110100001 : VALUE=19'b0000000_100001001010;
      15'b011_101110100010 : VALUE=19'b0000000_100001001010;
      15'b011_101110100011 : VALUE=19'b0000000_100001001010;
      15'b011_101110100100 : VALUE=19'b0000000_100001001010;
      15'b011_101110100101 : VALUE=19'b0000000_100001001001;
      15'b011_101110100110 : VALUE=19'b0000000_100001001001;
      15'b011_101110100111 : VALUE=19'b0000000_100001001001;
      15'b011_101110101000 : VALUE=19'b0000000_100001001001;
      15'b011_101110101001 : VALUE=19'b0000000_100001001001;
      15'b011_101110101010 : VALUE=19'b0000000_100001001001;
      15'b011_101110101011 : VALUE=19'b0000000_100001001001;
      15'b011_101110101100 : VALUE=19'b0000000_100001001001;
      15'b011_101110101101 : VALUE=19'b0000000_100001001001;
      15'b011_101110101110 : VALUE=19'b0000000_100001001001;
      15'b011_101110101111 : VALUE=19'b0000000_100001001001;
      15'b011_101110110000 : VALUE=19'b0000000_100001001001;
      15'b011_101110110001 : VALUE=19'b0000000_100001001001;
      15'b011_101110110010 : VALUE=19'b0000000_100001001001;
      15'b011_101110110011 : VALUE=19'b0000000_100001001000;
      15'b011_101110110100 : VALUE=19'b0000000_100001001000;
      15'b011_101110110101 : VALUE=19'b0000000_100001001000;
      15'b011_101110110110 : VALUE=19'b0000000_100001001000;
      15'b011_101110110111 : VALUE=19'b0000000_100001001000;
      15'b011_101110111000 : VALUE=19'b0000000_100001001000;
      15'b011_101110111001 : VALUE=19'b0000000_100001001000;
      15'b011_101110111010 : VALUE=19'b0000000_100001001000;
      15'b011_101110111011 : VALUE=19'b0000000_100001001000;
      15'b011_101110111100 : VALUE=19'b0000000_100001001000;
      15'b011_101110111101 : VALUE=19'b0000000_100001001000;
      15'b011_101110111110 : VALUE=19'b0000000_100001001000;
      15'b011_101110111111 : VALUE=19'b0000000_100001001000;
      15'b011_101111000000 : VALUE=19'b0000000_100001001000;
      15'b011_101111000001 : VALUE=19'b0000000_100001001000;
      15'b011_101111000010 : VALUE=19'b0000000_100001000111;
      15'b011_101111000011 : VALUE=19'b0000000_100001000111;
      15'b011_101111000100 : VALUE=19'b0000000_100001000111;
      15'b011_101111000101 : VALUE=19'b0000000_100001000111;
      15'b011_101111000110 : VALUE=19'b0000000_100001000111;
      15'b011_101111000111 : VALUE=19'b0000000_100001000111;
      15'b011_101111001000 : VALUE=19'b0000000_100001000111;
      15'b011_101111001001 : VALUE=19'b0000000_100001000111;
      15'b011_101111001010 : VALUE=19'b0000000_100001000111;
      15'b011_101111001011 : VALUE=19'b0000000_100001000111;
      15'b011_101111001100 : VALUE=19'b0000000_100001000111;
      15'b011_101111001101 : VALUE=19'b0000000_100001000111;
      15'b011_101111001110 : VALUE=19'b0000000_100001000111;
      15'b011_101111001111 : VALUE=19'b0000000_100001000111;
      15'b011_101111010000 : VALUE=19'b0000000_100001000110;
      15'b011_101111010001 : VALUE=19'b0000000_100001000110;
      15'b011_101111010010 : VALUE=19'b0000000_100001000110;
      15'b011_101111010011 : VALUE=19'b0000000_100001000110;
      15'b011_101111010100 : VALUE=19'b0000000_100001000110;
      15'b011_101111010101 : VALUE=19'b0000000_100001000110;
      15'b011_101111010110 : VALUE=19'b0000000_100001000110;
      15'b011_101111010111 : VALUE=19'b0000000_100001000110;
      15'b011_101111011000 : VALUE=19'b0000000_100001000110;
      15'b011_101111011001 : VALUE=19'b0000000_100001000110;
      15'b011_101111011010 : VALUE=19'b0000000_100001000110;
      15'b011_101111011011 : VALUE=19'b0000000_100001000110;
      15'b011_101111011100 : VALUE=19'b0000000_100001000110;
      15'b011_101111011101 : VALUE=19'b0000000_100001000110;
      15'b011_101111011110 : VALUE=19'b0000000_100001000110;
      15'b011_101111011111 : VALUE=19'b0000000_100001000101;
      15'b011_101111100000 : VALUE=19'b0000000_100001000101;
      15'b011_101111100001 : VALUE=19'b0000000_100001000101;
      15'b011_101111100010 : VALUE=19'b0000000_100001000101;
      15'b011_101111100011 : VALUE=19'b0000000_100001000101;
      15'b011_101111100100 : VALUE=19'b0000000_100001000101;
      15'b011_101111100101 : VALUE=19'b0000000_100001000101;
      15'b011_101111100110 : VALUE=19'b0000000_100001000101;
      15'b011_101111100111 : VALUE=19'b0000000_100001000101;
      15'b011_101111101000 : VALUE=19'b0000000_100001000101;
      15'b011_101111101001 : VALUE=19'b0000000_100001000101;
      15'b011_101111101010 : VALUE=19'b0000000_100001000101;
      15'b011_101111101011 : VALUE=19'b0000000_100001000101;
      15'b011_101111101100 : VALUE=19'b0000000_100001000101;
      15'b011_101111101101 : VALUE=19'b0000000_100001000100;
      15'b011_101111101110 : VALUE=19'b0000000_100001000100;
      15'b011_101111101111 : VALUE=19'b0000000_100001000100;
      15'b011_101111110000 : VALUE=19'b0000000_100001000100;
      15'b011_101111110001 : VALUE=19'b0000000_100001000100;
      15'b011_101111110010 : VALUE=19'b0000000_100001000100;
      15'b011_101111110011 : VALUE=19'b0000000_100001000100;
      15'b011_101111110100 : VALUE=19'b0000000_100001000100;
      15'b011_101111110101 : VALUE=19'b0000000_100001000100;
      15'b011_101111110110 : VALUE=19'b0000000_100001000100;
      15'b011_101111110111 : VALUE=19'b0000000_100001000100;
      15'b011_101111111000 : VALUE=19'b0000000_100001000100;
      15'b011_101111111001 : VALUE=19'b0000000_100001000100;
      15'b011_101111111010 : VALUE=19'b0000000_100001000100;
      15'b011_101111111011 : VALUE=19'b0000000_100001000100;
      15'b011_101111111100 : VALUE=19'b0000000_100001000011;
      15'b011_101111111101 : VALUE=19'b0000000_100001000011;
      15'b011_101111111110 : VALUE=19'b0000000_100001000011;
      15'b011_101111111111 : VALUE=19'b0000000_100001000011;
      15'b011_110000000000 : VALUE=19'b0000000_100001000011;
      15'b011_110000000001 : VALUE=19'b0000000_100001000011;
      15'b011_110000000010 : VALUE=19'b0000000_100001000011;
      15'b011_110000000011 : VALUE=19'b0000000_100001000011;
      15'b011_110000000100 : VALUE=19'b0000000_100001000011;
      15'b011_110000000101 : VALUE=19'b0000000_100001000011;
      15'b011_110000000110 : VALUE=19'b0000000_100001000011;
      15'b011_110000000111 : VALUE=19'b0000000_100001000011;
      15'b011_110000001000 : VALUE=19'b0000000_100001000011;
      15'b011_110000001001 : VALUE=19'b0000000_100001000011;
      15'b011_110000001010 : VALUE=19'b0000000_100001000010;
      15'b011_110000001011 : VALUE=19'b0000000_100001000010;
      15'b011_110000001100 : VALUE=19'b0000000_100001000010;
      15'b011_110000001101 : VALUE=19'b0000000_100001000010;
      15'b011_110000001110 : VALUE=19'b0000000_100001000010;
      15'b011_110000001111 : VALUE=19'b0000000_100001000010;
      15'b011_110000010000 : VALUE=19'b0000000_100001000010;
      15'b011_110000010001 : VALUE=19'b0000000_100001000010;
      15'b011_110000010010 : VALUE=19'b0000000_100001000010;
      15'b011_110000010011 : VALUE=19'b0000000_100001000010;
      15'b011_110000010100 : VALUE=19'b0000000_100001000010;
      15'b011_110000010101 : VALUE=19'b0000000_100001000010;
      15'b011_110000010110 : VALUE=19'b0000000_100001000010;
      15'b011_110000010111 : VALUE=19'b0000000_100001000010;
      15'b011_110000011000 : VALUE=19'b0000000_100001000010;
      15'b011_110000011001 : VALUE=19'b0000000_100001000001;
      15'b011_110000011010 : VALUE=19'b0000000_100001000001;
      15'b011_110000011011 : VALUE=19'b0000000_100001000001;
      15'b011_110000011100 : VALUE=19'b0000000_100001000001;
      15'b011_110000011101 : VALUE=19'b0000000_100001000001;
      15'b011_110000011110 : VALUE=19'b0000000_100001000001;
      15'b011_110000011111 : VALUE=19'b0000000_100001000001;
      15'b011_110000100000 : VALUE=19'b0000000_100001000001;
      15'b011_110000100001 : VALUE=19'b0000000_100001000001;
      15'b011_110000100010 : VALUE=19'b0000000_100001000001;
      15'b011_110000100011 : VALUE=19'b0000000_100001000001;
      15'b011_110000100100 : VALUE=19'b0000000_100001000001;
      15'b011_110000100101 : VALUE=19'b0000000_100001000001;
      15'b011_110000100110 : VALUE=19'b0000000_100001000001;
      15'b011_110000100111 : VALUE=19'b0000000_100001000000;
      15'b011_110000101000 : VALUE=19'b0000000_100001000000;
      15'b011_110000101001 : VALUE=19'b0000000_100001000000;
      15'b011_110000101010 : VALUE=19'b0000000_100001000000;
      15'b011_110000101011 : VALUE=19'b0000000_100001000000;
      15'b011_110000101100 : VALUE=19'b0000000_100001000000;
      15'b011_110000101101 : VALUE=19'b0000000_100001000000;
      15'b011_110000101110 : VALUE=19'b0000000_100001000000;
      15'b011_110000101111 : VALUE=19'b0000000_100001000000;
      15'b011_110000110000 : VALUE=19'b0000000_100001000000;
      15'b011_110000110001 : VALUE=19'b0000000_100001000000;
      15'b011_110000110010 : VALUE=19'b0000000_100001000000;
      15'b011_110000110011 : VALUE=19'b0000000_100001000000;
      15'b011_110000110100 : VALUE=19'b0000000_100001000000;
      15'b011_110000110101 : VALUE=19'b0000000_100001000000;
      15'b011_110000110110 : VALUE=19'b0000000_100000111111;
      15'b011_110000110111 : VALUE=19'b0000000_100000111111;
      15'b011_110000111000 : VALUE=19'b0000000_100000111111;
      15'b011_110000111001 : VALUE=19'b0000000_100000111111;
      15'b011_110000111010 : VALUE=19'b0000000_100000111111;
      15'b011_110000111011 : VALUE=19'b0000000_100000111111;
      15'b011_110000111100 : VALUE=19'b0000000_100000111111;
      15'b011_110000111101 : VALUE=19'b0000000_100000111111;
      15'b011_110000111110 : VALUE=19'b0000000_100000111111;
      15'b011_110000111111 : VALUE=19'b0000000_100000111111;
      15'b011_110001000000 : VALUE=19'b0000000_100000111111;
      15'b011_110001000001 : VALUE=19'b0000000_100000111111;
      15'b011_110001000010 : VALUE=19'b0000000_100000111111;
      15'b011_110001000011 : VALUE=19'b0000000_100000111111;
      15'b011_110001000100 : VALUE=19'b0000000_100000111110;
      15'b011_110001000101 : VALUE=19'b0000000_100000111110;
      15'b011_110001000110 : VALUE=19'b0000000_100000111110;
      15'b011_110001000111 : VALUE=19'b0000000_100000111110;
      15'b011_110001001000 : VALUE=19'b0000000_100000111110;
      15'b011_110001001001 : VALUE=19'b0000000_100000111110;
      15'b011_110001001010 : VALUE=19'b0000000_100000111110;
      15'b011_110001001011 : VALUE=19'b0000000_100000111110;
      15'b011_110001001100 : VALUE=19'b0000000_100000111110;
      15'b011_110001001101 : VALUE=19'b0000000_100000111110;
      15'b011_110001001110 : VALUE=19'b0000000_100000111110;
      15'b011_110001001111 : VALUE=19'b0000000_100000111110;
      15'b011_110001010000 : VALUE=19'b0000000_100000111110;
      15'b011_110001010001 : VALUE=19'b0000000_100000111110;
      15'b011_110001010010 : VALUE=19'b0000000_100000111110;
      15'b011_110001010011 : VALUE=19'b0000000_100000111101;
      15'b011_110001010100 : VALUE=19'b0000000_100000111101;
      15'b011_110001010101 : VALUE=19'b0000000_100000111101;
      15'b011_110001010110 : VALUE=19'b0000000_100000111101;
      15'b011_110001010111 : VALUE=19'b0000000_100000111101;
      15'b011_110001011000 : VALUE=19'b0000000_100000111101;
      15'b011_110001011001 : VALUE=19'b0000000_100000111101;
      15'b011_110001011010 : VALUE=19'b0000000_100000111101;
      15'b011_110001011011 : VALUE=19'b0000000_100000111101;
      15'b011_110001011100 : VALUE=19'b0000000_100000111101;
      15'b011_110001011101 : VALUE=19'b0000000_100000111101;
      15'b011_110001011110 : VALUE=19'b0000000_100000111101;
      15'b011_110001011111 : VALUE=19'b0000000_100000111101;
      15'b011_110001100000 : VALUE=19'b0000000_100000111101;
      15'b011_110001100001 : VALUE=19'b0000000_100000111101;
      15'b011_110001100010 : VALUE=19'b0000000_100000111100;
      15'b011_110001100011 : VALUE=19'b0000000_100000111100;
      15'b011_110001100100 : VALUE=19'b0000000_100000111100;
      15'b011_110001100101 : VALUE=19'b0000000_100000111100;
      15'b011_110001100110 : VALUE=19'b0000000_100000111100;
      15'b011_110001100111 : VALUE=19'b0000000_100000111100;
      15'b011_110001101000 : VALUE=19'b0000000_100000111100;
      15'b011_110001101001 : VALUE=19'b0000000_100000111100;
      15'b011_110001101010 : VALUE=19'b0000000_100000111100;
      15'b011_110001101011 : VALUE=19'b0000000_100000111100;
      15'b011_110001101100 : VALUE=19'b0000000_100000111100;
      15'b011_110001101101 : VALUE=19'b0000000_100000111100;
      15'b011_110001101110 : VALUE=19'b0000000_100000111100;
      15'b011_110001101111 : VALUE=19'b0000000_100000111100;
      15'b011_110001110000 : VALUE=19'b0000000_100000111011;
      15'b011_110001110001 : VALUE=19'b0000000_100000111011;
      15'b011_110001110010 : VALUE=19'b0000000_100000111011;
      15'b011_110001110011 : VALUE=19'b0000000_100000111011;
      15'b011_110001110100 : VALUE=19'b0000000_100000111011;
      15'b011_110001110101 : VALUE=19'b0000000_100000111011;
      15'b011_110001110110 : VALUE=19'b0000000_100000111011;
      15'b011_110001110111 : VALUE=19'b0000000_100000111011;
      15'b011_110001111000 : VALUE=19'b0000000_100000111011;
      15'b011_110001111001 : VALUE=19'b0000000_100000111011;
      15'b011_110001111010 : VALUE=19'b0000000_100000111011;
      15'b011_110001111011 : VALUE=19'b0000000_100000111011;
      15'b011_110001111100 : VALUE=19'b0000000_100000111011;
      15'b011_110001111101 : VALUE=19'b0000000_100000111011;
      15'b011_110001111110 : VALUE=19'b0000000_100000111011;
      15'b011_110001111111 : VALUE=19'b0000000_100000111010;
      15'b011_110010000000 : VALUE=19'b0000000_100000111010;
      15'b011_110010000001 : VALUE=19'b0000000_100000111010;
      15'b011_110010000010 : VALUE=19'b0000000_100000111010;
      15'b011_110010000011 : VALUE=19'b0000000_100000111010;
      15'b011_110010000100 : VALUE=19'b0000000_100000111010;
      15'b011_110010000101 : VALUE=19'b0000000_100000111010;
      15'b011_110010000110 : VALUE=19'b0000000_100000111010;
      15'b011_110010000111 : VALUE=19'b0000000_100000111010;
      15'b011_110010001000 : VALUE=19'b0000000_100000111010;
      15'b011_110010001001 : VALUE=19'b0000000_100000111010;
      15'b011_110010001010 : VALUE=19'b0000000_100000111010;
      15'b011_110010001011 : VALUE=19'b0000000_100000111010;
      15'b011_110010001100 : VALUE=19'b0000000_100000111010;
      15'b011_110010001101 : VALUE=19'b0000000_100000111010;
      15'b011_110010001110 : VALUE=19'b0000000_100000111001;
      15'b011_110010001111 : VALUE=19'b0000000_100000111001;
      15'b011_110010010000 : VALUE=19'b0000000_100000111001;
      15'b011_110010010001 : VALUE=19'b0000000_100000111001;
      15'b011_110010010010 : VALUE=19'b0000000_100000111001;
      15'b011_110010010011 : VALUE=19'b0000000_100000111001;
      15'b011_110010010100 : VALUE=19'b0000000_100000111001;
      15'b011_110010010101 : VALUE=19'b0000000_100000111001;
      15'b011_110010010110 : VALUE=19'b0000000_100000111001;
      15'b011_110010010111 : VALUE=19'b0000000_100000111001;
      15'b011_110010011000 : VALUE=19'b0000000_100000111001;
      15'b011_110010011001 : VALUE=19'b0000000_100000111001;
      15'b011_110010011010 : VALUE=19'b0000000_100000111001;
      15'b011_110010011011 : VALUE=19'b0000000_100000111001;
      15'b011_110010011100 : VALUE=19'b0000000_100000111001;
      15'b011_110010011101 : VALUE=19'b0000000_100000111000;
      15'b011_110010011110 : VALUE=19'b0000000_100000111000;
      15'b011_110010011111 : VALUE=19'b0000000_100000111000;
      15'b011_110010100000 : VALUE=19'b0000000_100000111000;
      15'b011_110010100001 : VALUE=19'b0000000_100000111000;
      15'b011_110010100010 : VALUE=19'b0000000_100000111000;
      15'b011_110010100011 : VALUE=19'b0000000_100000111000;
      15'b011_110010100100 : VALUE=19'b0000000_100000111000;
      15'b011_110010100101 : VALUE=19'b0000000_100000111000;
      15'b011_110010100110 : VALUE=19'b0000000_100000111000;
      15'b011_110010100111 : VALUE=19'b0000000_100000111000;
      15'b011_110010101000 : VALUE=19'b0000000_100000111000;
      15'b011_110010101001 : VALUE=19'b0000000_100000111000;
      15'b011_110010101010 : VALUE=19'b0000000_100000111000;
      15'b011_110010101011 : VALUE=19'b0000000_100000110111;
      15'b011_110010101100 : VALUE=19'b0000000_100000110111;
      15'b011_110010101101 : VALUE=19'b0000000_100000110111;
      15'b011_110010101110 : VALUE=19'b0000000_100000110111;
      15'b011_110010101111 : VALUE=19'b0000000_100000110111;
      15'b011_110010110000 : VALUE=19'b0000000_100000110111;
      15'b011_110010110001 : VALUE=19'b0000000_100000110111;
      15'b011_110010110010 : VALUE=19'b0000000_100000110111;
      15'b011_110010110011 : VALUE=19'b0000000_100000110111;
      15'b011_110010110100 : VALUE=19'b0000000_100000110111;
      15'b011_110010110101 : VALUE=19'b0000000_100000110111;
      15'b011_110010110110 : VALUE=19'b0000000_100000110111;
      15'b011_110010110111 : VALUE=19'b0000000_100000110111;
      15'b011_110010111000 : VALUE=19'b0000000_100000110111;
      15'b011_110010111001 : VALUE=19'b0000000_100000110111;
      15'b011_110010111010 : VALUE=19'b0000000_100000110110;
      15'b011_110010111011 : VALUE=19'b0000000_100000110110;
      15'b011_110010111100 : VALUE=19'b0000000_100000110110;
      15'b011_110010111101 : VALUE=19'b0000000_100000110110;
      15'b011_110010111110 : VALUE=19'b0000000_100000110110;
      15'b011_110010111111 : VALUE=19'b0000000_100000110110;
      15'b011_110011000000 : VALUE=19'b0000000_100000110110;
      15'b011_110011000001 : VALUE=19'b0000000_100000110110;
      15'b011_110011000010 : VALUE=19'b0000000_100000110110;
      15'b011_110011000011 : VALUE=19'b0000000_100000110110;
      15'b011_110011000100 : VALUE=19'b0000000_100000110110;
      15'b011_110011000101 : VALUE=19'b0000000_100000110110;
      15'b011_110011000110 : VALUE=19'b0000000_100000110110;
      15'b011_110011000111 : VALUE=19'b0000000_100000110110;
      15'b011_110011001000 : VALUE=19'b0000000_100000110110;
      15'b011_110011001001 : VALUE=19'b0000000_100000110101;
      15'b011_110011001010 : VALUE=19'b0000000_100000110101;
      15'b011_110011001011 : VALUE=19'b0000000_100000110101;
      15'b011_110011001100 : VALUE=19'b0000000_100000110101;
      15'b011_110011001101 : VALUE=19'b0000000_100000110101;
      15'b011_110011001110 : VALUE=19'b0000000_100000110101;
      15'b011_110011001111 : VALUE=19'b0000000_100000110101;
      15'b011_110011010000 : VALUE=19'b0000000_100000110101;
      15'b011_110011010001 : VALUE=19'b0000000_100000110101;
      15'b011_110011010010 : VALUE=19'b0000000_100000110101;
      15'b011_110011010011 : VALUE=19'b0000000_100000110101;
      15'b011_110011010100 : VALUE=19'b0000000_100000110101;
      15'b011_110011010101 : VALUE=19'b0000000_100000110101;
      15'b011_110011010110 : VALUE=19'b0000000_100000110101;
      15'b011_110011010111 : VALUE=19'b0000000_100000110101;
      15'b011_110011011000 : VALUE=19'b0000000_100000110100;
      15'b011_110011011001 : VALUE=19'b0000000_100000110100;
      15'b011_110011011010 : VALUE=19'b0000000_100000110100;
      15'b011_110011011011 : VALUE=19'b0000000_100000110100;
      15'b011_110011011100 : VALUE=19'b0000000_100000110100;
      15'b011_110011011101 : VALUE=19'b0000000_100000110100;
      15'b011_110011011110 : VALUE=19'b0000000_100000110100;
      15'b011_110011011111 : VALUE=19'b0000000_100000110100;
      15'b011_110011100000 : VALUE=19'b0000000_100000110100;
      15'b011_110011100001 : VALUE=19'b0000000_100000110100;
      15'b011_110011100010 : VALUE=19'b0000000_100000110100;
      15'b011_110011100011 : VALUE=19'b0000000_100000110100;
      15'b011_110011100100 : VALUE=19'b0000000_100000110100;
      15'b011_110011100101 : VALUE=19'b0000000_100000110100;
      15'b011_110011100110 : VALUE=19'b0000000_100000110100;
      15'b011_110011100111 : VALUE=19'b0000000_100000110011;
      15'b011_110011101000 : VALUE=19'b0000000_100000110011;
      15'b011_110011101001 : VALUE=19'b0000000_100000110011;
      15'b011_110011101010 : VALUE=19'b0000000_100000110011;
      15'b011_110011101011 : VALUE=19'b0000000_100000110011;
      15'b011_110011101100 : VALUE=19'b0000000_100000110011;
      15'b011_110011101101 : VALUE=19'b0000000_100000110011;
      15'b011_110011101110 : VALUE=19'b0000000_100000110011;
      15'b011_110011101111 : VALUE=19'b0000000_100000110011;
      15'b011_110011110000 : VALUE=19'b0000000_100000110011;
      15'b011_110011110001 : VALUE=19'b0000000_100000110011;
      15'b011_110011110010 : VALUE=19'b0000000_100000110011;
      15'b011_110011110011 : VALUE=19'b0000000_100000110011;
      15'b011_110011110100 : VALUE=19'b0000000_100000110011;
      15'b011_110011110101 : VALUE=19'b0000000_100000110010;
      15'b011_110011110110 : VALUE=19'b0000000_100000110010;
      15'b011_110011110111 : VALUE=19'b0000000_100000110010;
      15'b011_110011111000 : VALUE=19'b0000000_100000110010;
      15'b011_110011111001 : VALUE=19'b0000000_100000110010;
      15'b011_110011111010 : VALUE=19'b0000000_100000110010;
      15'b011_110011111011 : VALUE=19'b0000000_100000110010;
      15'b011_110011111100 : VALUE=19'b0000000_100000110010;
      15'b011_110011111101 : VALUE=19'b0000000_100000110010;
      15'b011_110011111110 : VALUE=19'b0000000_100000110010;
      15'b011_110011111111 : VALUE=19'b0000000_100000110010;
      15'b011_110100000000 : VALUE=19'b0000000_100000110010;
      15'b011_110100000001 : VALUE=19'b0000000_100000110010;
      15'b011_110100000010 : VALUE=19'b0000000_100000110010;
      15'b011_110100000011 : VALUE=19'b0000000_100000110010;
      15'b011_110100000100 : VALUE=19'b0000000_100000110001;
      15'b011_110100000101 : VALUE=19'b0000000_100000110001;
      15'b011_110100000110 : VALUE=19'b0000000_100000110001;
      15'b011_110100000111 : VALUE=19'b0000000_100000110001;
      15'b011_110100001000 : VALUE=19'b0000000_100000110001;
      15'b011_110100001001 : VALUE=19'b0000000_100000110001;
      15'b011_110100001010 : VALUE=19'b0000000_100000110001;
      15'b011_110100001011 : VALUE=19'b0000000_100000110001;
      15'b011_110100001100 : VALUE=19'b0000000_100000110001;
      15'b011_110100001101 : VALUE=19'b0000000_100000110001;
      15'b011_110100001110 : VALUE=19'b0000000_100000110001;
      15'b011_110100001111 : VALUE=19'b0000000_100000110001;
      15'b011_110100010000 : VALUE=19'b0000000_100000110001;
      15'b011_110100010001 : VALUE=19'b0000000_100000110001;
      15'b011_110100010010 : VALUE=19'b0000000_100000110001;
      15'b011_110100010011 : VALUE=19'b0000000_100000110000;
      15'b011_110100010100 : VALUE=19'b0000000_100000110000;
      15'b011_110100010101 : VALUE=19'b0000000_100000110000;
      15'b011_110100010110 : VALUE=19'b0000000_100000110000;
      15'b011_110100010111 : VALUE=19'b0000000_100000110000;
      15'b011_110100011000 : VALUE=19'b0000000_100000110000;
      15'b011_110100011001 : VALUE=19'b0000000_100000110000;
      15'b011_110100011010 : VALUE=19'b0000000_100000110000;
      15'b011_110100011011 : VALUE=19'b0000000_100000110000;
      15'b011_110100011100 : VALUE=19'b0000000_100000110000;
      15'b011_110100011101 : VALUE=19'b0000000_100000110000;
      15'b011_110100011110 : VALUE=19'b0000000_100000110000;
      15'b011_110100011111 : VALUE=19'b0000000_100000110000;
      15'b011_110100100000 : VALUE=19'b0000000_100000110000;
      15'b011_110100100001 : VALUE=19'b0000000_100000110000;
      15'b011_110100100010 : VALUE=19'b0000000_100000101111;
      15'b011_110100100011 : VALUE=19'b0000000_100000101111;
      15'b011_110100100100 : VALUE=19'b0000000_100000101111;
      15'b011_110100100101 : VALUE=19'b0000000_100000101111;
      15'b011_110100100110 : VALUE=19'b0000000_100000101111;
      15'b011_110100100111 : VALUE=19'b0000000_100000101111;
      15'b011_110100101000 : VALUE=19'b0000000_100000101111;
      15'b011_110100101001 : VALUE=19'b0000000_100000101111;
      15'b011_110100101010 : VALUE=19'b0000000_100000101111;
      15'b011_110100101011 : VALUE=19'b0000000_100000101111;
      15'b011_110100101100 : VALUE=19'b0000000_100000101111;
      15'b011_110100101101 : VALUE=19'b0000000_100000101111;
      15'b011_110100101110 : VALUE=19'b0000000_100000101111;
      15'b011_110100101111 : VALUE=19'b0000000_100000101111;
      15'b011_110100110000 : VALUE=19'b0000000_100000101111;
      15'b011_110100110001 : VALUE=19'b0000000_100000101110;
      15'b011_110100110010 : VALUE=19'b0000000_100000101110;
      15'b011_110100110011 : VALUE=19'b0000000_100000101110;
      15'b011_110100110100 : VALUE=19'b0000000_100000101110;
      15'b011_110100110101 : VALUE=19'b0000000_100000101110;
      15'b011_110100110110 : VALUE=19'b0000000_100000101110;
      15'b011_110100110111 : VALUE=19'b0000000_100000101110;
      15'b011_110100111000 : VALUE=19'b0000000_100000101110;
      15'b011_110100111001 : VALUE=19'b0000000_100000101110;
      15'b011_110100111010 : VALUE=19'b0000000_100000101110;
      15'b011_110100111011 : VALUE=19'b0000000_100000101110;
      15'b011_110100111100 : VALUE=19'b0000000_100000101110;
      15'b011_110100111101 : VALUE=19'b0000000_100000101110;
      15'b011_110100111110 : VALUE=19'b0000000_100000101110;
      15'b011_110100111111 : VALUE=19'b0000000_100000101110;
      15'b011_110101000000 : VALUE=19'b0000000_100000101101;
      15'b011_110101000001 : VALUE=19'b0000000_100000101101;
      15'b011_110101000010 : VALUE=19'b0000000_100000101101;
      15'b011_110101000011 : VALUE=19'b0000000_100000101101;
      15'b011_110101000100 : VALUE=19'b0000000_100000101101;
      15'b011_110101000101 : VALUE=19'b0000000_100000101101;
      15'b011_110101000110 : VALUE=19'b0000000_100000101101;
      15'b011_110101000111 : VALUE=19'b0000000_100000101101;
      15'b011_110101001000 : VALUE=19'b0000000_100000101101;
      15'b011_110101001001 : VALUE=19'b0000000_100000101101;
      15'b011_110101001010 : VALUE=19'b0000000_100000101101;
      15'b011_110101001011 : VALUE=19'b0000000_100000101101;
      15'b011_110101001100 : VALUE=19'b0000000_100000101101;
      15'b011_110101001101 : VALUE=19'b0000000_100000101101;
      15'b011_110101001110 : VALUE=19'b0000000_100000101101;
      15'b011_110101001111 : VALUE=19'b0000000_100000101100;
      15'b011_110101010000 : VALUE=19'b0000000_100000101100;
      15'b011_110101010001 : VALUE=19'b0000000_100000101100;
      15'b011_110101010010 : VALUE=19'b0000000_100000101100;
      15'b011_110101010011 : VALUE=19'b0000000_100000101100;
      15'b011_110101010100 : VALUE=19'b0000000_100000101100;
      15'b011_110101010101 : VALUE=19'b0000000_100000101100;
      15'b011_110101010110 : VALUE=19'b0000000_100000101100;
      15'b011_110101010111 : VALUE=19'b0000000_100000101100;
      15'b011_110101011000 : VALUE=19'b0000000_100000101100;
      15'b011_110101011001 : VALUE=19'b0000000_100000101100;
      15'b011_110101011010 : VALUE=19'b0000000_100000101100;
      15'b011_110101011011 : VALUE=19'b0000000_100000101100;
      15'b011_110101011100 : VALUE=19'b0000000_100000101100;
      15'b011_110101011101 : VALUE=19'b0000000_100000101100;
      15'b011_110101011110 : VALUE=19'b0000000_100000101011;
      15'b011_110101011111 : VALUE=19'b0000000_100000101011;
      15'b011_110101100000 : VALUE=19'b0000000_100000101011;
      15'b011_110101100001 : VALUE=19'b0000000_100000101011;
      15'b011_110101100010 : VALUE=19'b0000000_100000101011;
      15'b011_110101100011 : VALUE=19'b0000000_100000101011;
      15'b011_110101100100 : VALUE=19'b0000000_100000101011;
      15'b011_110101100101 : VALUE=19'b0000000_100000101011;
      15'b011_110101100110 : VALUE=19'b0000000_100000101011;
      15'b011_110101100111 : VALUE=19'b0000000_100000101011;
      15'b011_110101101000 : VALUE=19'b0000000_100000101011;
      15'b011_110101101001 : VALUE=19'b0000000_100000101011;
      15'b011_110101101010 : VALUE=19'b0000000_100000101011;
      15'b011_110101101011 : VALUE=19'b0000000_100000101011;
      15'b011_110101101100 : VALUE=19'b0000000_100000101011;
      15'b011_110101101101 : VALUE=19'b0000000_100000101010;
      15'b011_110101101110 : VALUE=19'b0000000_100000101010;
      15'b011_110101101111 : VALUE=19'b0000000_100000101010;
      15'b011_110101110000 : VALUE=19'b0000000_100000101010;
      15'b011_110101110001 : VALUE=19'b0000000_100000101010;
      15'b011_110101110010 : VALUE=19'b0000000_100000101010;
      15'b011_110101110011 : VALUE=19'b0000000_100000101010;
      15'b011_110101110100 : VALUE=19'b0000000_100000101010;
      15'b011_110101110101 : VALUE=19'b0000000_100000101010;
      15'b011_110101110110 : VALUE=19'b0000000_100000101010;
      15'b011_110101110111 : VALUE=19'b0000000_100000101010;
      15'b011_110101111000 : VALUE=19'b0000000_100000101010;
      15'b011_110101111001 : VALUE=19'b0000000_100000101010;
      15'b011_110101111010 : VALUE=19'b0000000_100000101010;
      15'b011_110101111011 : VALUE=19'b0000000_100000101010;
      15'b011_110101111100 : VALUE=19'b0000000_100000101001;
      15'b011_110101111101 : VALUE=19'b0000000_100000101001;
      15'b011_110101111110 : VALUE=19'b0000000_100000101001;
      15'b011_110101111111 : VALUE=19'b0000000_100000101001;
      15'b011_110110000000 : VALUE=19'b0000000_100000101001;
      15'b011_110110000001 : VALUE=19'b0000000_100000101001;
      15'b011_110110000010 : VALUE=19'b0000000_100000101001;
      15'b011_110110000011 : VALUE=19'b0000000_100000101001;
      15'b011_110110000100 : VALUE=19'b0000000_100000101001;
      15'b011_110110000101 : VALUE=19'b0000000_100000101001;
      15'b011_110110000110 : VALUE=19'b0000000_100000101001;
      15'b011_110110000111 : VALUE=19'b0000000_100000101001;
      15'b011_110110001000 : VALUE=19'b0000000_100000101001;
      15'b011_110110001001 : VALUE=19'b0000000_100000101001;
      15'b011_110110001010 : VALUE=19'b0000000_100000101001;
      15'b011_110110001011 : VALUE=19'b0000000_100000101000;
      15'b011_110110001100 : VALUE=19'b0000000_100000101000;
      15'b011_110110001101 : VALUE=19'b0000000_100000101000;
      15'b011_110110001110 : VALUE=19'b0000000_100000101000;
      15'b011_110110001111 : VALUE=19'b0000000_100000101000;
      15'b011_110110010000 : VALUE=19'b0000000_100000101000;
      15'b011_110110010001 : VALUE=19'b0000000_100000101000;
      15'b011_110110010010 : VALUE=19'b0000000_100000101000;
      15'b011_110110010011 : VALUE=19'b0000000_100000101000;
      15'b011_110110010100 : VALUE=19'b0000000_100000101000;
      15'b011_110110010101 : VALUE=19'b0000000_100000101000;
      15'b011_110110010110 : VALUE=19'b0000000_100000101000;
      15'b011_110110010111 : VALUE=19'b0000000_100000101000;
      15'b011_110110011000 : VALUE=19'b0000000_100000101000;
      15'b011_110110011001 : VALUE=19'b0000000_100000101000;
      15'b011_110110011010 : VALUE=19'b0000000_100000100111;
      15'b011_110110011011 : VALUE=19'b0000000_100000100111;
      15'b011_110110011100 : VALUE=19'b0000000_100000100111;
      15'b011_110110011101 : VALUE=19'b0000000_100000100111;
      15'b011_110110011110 : VALUE=19'b0000000_100000100111;
      15'b011_110110011111 : VALUE=19'b0000000_100000100111;
      15'b011_110110100000 : VALUE=19'b0000000_100000100111;
      15'b011_110110100001 : VALUE=19'b0000000_100000100111;
      15'b011_110110100010 : VALUE=19'b0000000_100000100111;
      15'b011_110110100011 : VALUE=19'b0000000_100000100111;
      15'b011_110110100100 : VALUE=19'b0000000_100000100111;
      15'b011_110110100101 : VALUE=19'b0000000_100000100111;
      15'b011_110110100110 : VALUE=19'b0000000_100000100111;
      15'b011_110110100111 : VALUE=19'b0000000_100000100111;
      15'b011_110110101000 : VALUE=19'b0000000_100000100111;
      15'b011_110110101001 : VALUE=19'b0000000_100000100110;
      15'b011_110110101010 : VALUE=19'b0000000_100000100110;
      15'b011_110110101011 : VALUE=19'b0000000_100000100110;
      15'b011_110110101100 : VALUE=19'b0000000_100000100110;
      15'b011_110110101101 : VALUE=19'b0000000_100000100110;
      15'b011_110110101110 : VALUE=19'b0000000_100000100110;
      15'b011_110110101111 : VALUE=19'b0000000_100000100110;
      15'b011_110110110000 : VALUE=19'b0000000_100000100110;
      15'b011_110110110001 : VALUE=19'b0000000_100000100110;
      15'b011_110110110010 : VALUE=19'b0000000_100000100110;
      15'b011_110110110011 : VALUE=19'b0000000_100000100110;
      15'b011_110110110100 : VALUE=19'b0000000_100000100110;
      15'b011_110110110101 : VALUE=19'b0000000_100000100110;
      15'b011_110110110110 : VALUE=19'b0000000_100000100110;
      15'b011_110110110111 : VALUE=19'b0000000_100000100110;
      15'b011_110110111000 : VALUE=19'b0000000_100000100110;
      15'b011_110110111001 : VALUE=19'b0000000_100000100101;
      15'b011_110110111010 : VALUE=19'b0000000_100000100101;
      15'b011_110110111011 : VALUE=19'b0000000_100000100101;
      15'b011_110110111100 : VALUE=19'b0000000_100000100101;
      15'b011_110110111101 : VALUE=19'b0000000_100000100101;
      15'b011_110110111110 : VALUE=19'b0000000_100000100101;
      15'b011_110110111111 : VALUE=19'b0000000_100000100101;
      15'b011_110111000000 : VALUE=19'b0000000_100000100101;
      15'b011_110111000001 : VALUE=19'b0000000_100000100101;
      15'b011_110111000010 : VALUE=19'b0000000_100000100101;
      15'b011_110111000011 : VALUE=19'b0000000_100000100101;
      15'b011_110111000100 : VALUE=19'b0000000_100000100101;
      15'b011_110111000101 : VALUE=19'b0000000_100000100101;
      15'b011_110111000110 : VALUE=19'b0000000_100000100101;
      15'b011_110111000111 : VALUE=19'b0000000_100000100101;
      15'b011_110111001000 : VALUE=19'b0000000_100000100100;
      15'b011_110111001001 : VALUE=19'b0000000_100000100100;
      15'b011_110111001010 : VALUE=19'b0000000_100000100100;
      15'b011_110111001011 : VALUE=19'b0000000_100000100100;
      15'b011_110111001100 : VALUE=19'b0000000_100000100100;
      15'b011_110111001101 : VALUE=19'b0000000_100000100100;
      15'b011_110111001110 : VALUE=19'b0000000_100000100100;
      15'b011_110111001111 : VALUE=19'b0000000_100000100100;
      15'b011_110111010000 : VALUE=19'b0000000_100000100100;
      15'b011_110111010001 : VALUE=19'b0000000_100000100100;
      15'b011_110111010010 : VALUE=19'b0000000_100000100100;
      15'b011_110111010011 : VALUE=19'b0000000_100000100100;
      15'b011_110111010100 : VALUE=19'b0000000_100000100100;
      15'b011_110111010101 : VALUE=19'b0000000_100000100100;
      15'b011_110111010110 : VALUE=19'b0000000_100000100100;
      15'b011_110111010111 : VALUE=19'b0000000_100000100011;
      15'b011_110111011000 : VALUE=19'b0000000_100000100011;
      15'b011_110111011001 : VALUE=19'b0000000_100000100011;
      15'b011_110111011010 : VALUE=19'b0000000_100000100011;
      15'b011_110111011011 : VALUE=19'b0000000_100000100011;
      15'b011_110111011100 : VALUE=19'b0000000_100000100011;
      15'b011_110111011101 : VALUE=19'b0000000_100000100011;
      15'b011_110111011110 : VALUE=19'b0000000_100000100011;
      15'b011_110111011111 : VALUE=19'b0000000_100000100011;
      15'b011_110111100000 : VALUE=19'b0000000_100000100011;
      15'b011_110111100001 : VALUE=19'b0000000_100000100011;
      15'b011_110111100010 : VALUE=19'b0000000_100000100011;
      15'b011_110111100011 : VALUE=19'b0000000_100000100011;
      15'b011_110111100100 : VALUE=19'b0000000_100000100011;
      15'b011_110111100101 : VALUE=19'b0000000_100000100011;
      15'b011_110111100110 : VALUE=19'b0000000_100000100010;
      15'b011_110111100111 : VALUE=19'b0000000_100000100010;
      15'b011_110111101000 : VALUE=19'b0000000_100000100010;
      15'b011_110111101001 : VALUE=19'b0000000_100000100010;
      15'b011_110111101010 : VALUE=19'b0000000_100000100010;
      15'b011_110111101011 : VALUE=19'b0000000_100000100010;
      15'b011_110111101100 : VALUE=19'b0000000_100000100010;
      15'b011_110111101101 : VALUE=19'b0000000_100000100010;
      15'b011_110111101110 : VALUE=19'b0000000_100000100010;
      15'b011_110111101111 : VALUE=19'b0000000_100000100010;
      15'b011_110111110000 : VALUE=19'b0000000_100000100010;
      15'b011_110111110001 : VALUE=19'b0000000_100000100010;
      15'b011_110111110010 : VALUE=19'b0000000_100000100010;
      15'b011_110111110011 : VALUE=19'b0000000_100000100010;
      15'b011_110111110100 : VALUE=19'b0000000_100000100010;
      15'b011_110111110101 : VALUE=19'b0000000_100000100001;
      15'b011_110111110110 : VALUE=19'b0000000_100000100001;
      15'b011_110111110111 : VALUE=19'b0000000_100000100001;
      15'b011_110111111000 : VALUE=19'b0000000_100000100001;
      15'b011_110111111001 : VALUE=19'b0000000_100000100001;
      15'b011_110111111010 : VALUE=19'b0000000_100000100001;
      15'b011_110111111011 : VALUE=19'b0000000_100000100001;
      15'b011_110111111100 : VALUE=19'b0000000_100000100001;
      15'b011_110111111101 : VALUE=19'b0000000_100000100001;
      15'b011_110111111110 : VALUE=19'b0000000_100000100001;
      15'b011_110111111111 : VALUE=19'b0000000_100000100001;
      15'b011_111000000000 : VALUE=19'b0000000_100000100001;
      15'b011_111000000001 : VALUE=19'b0000000_100000100001;
      15'b011_111000000010 : VALUE=19'b0000000_100000100001;
      15'b011_111000000011 : VALUE=19'b0000000_100000100001;
      15'b011_111000000100 : VALUE=19'b0000000_100000100001;
      15'b011_111000000101 : VALUE=19'b0000000_100000100000;
      15'b011_111000000110 : VALUE=19'b0000000_100000100000;
      15'b011_111000000111 : VALUE=19'b0000000_100000100000;
      15'b011_111000001000 : VALUE=19'b0000000_100000100000;
      15'b011_111000001001 : VALUE=19'b0000000_100000100000;
      15'b011_111000001010 : VALUE=19'b0000000_100000100000;
      15'b011_111000001011 : VALUE=19'b0000000_100000100000;
      15'b011_111000001100 : VALUE=19'b0000000_100000100000;
      15'b011_111000001101 : VALUE=19'b0000000_100000100000;
      15'b011_111000001110 : VALUE=19'b0000000_100000100000;
      15'b011_111000001111 : VALUE=19'b0000000_100000100000;
      15'b011_111000010000 : VALUE=19'b0000000_100000100000;
      15'b011_111000010001 : VALUE=19'b0000000_100000100000;
      15'b011_111000010010 : VALUE=19'b0000000_100000100000;
      15'b011_111000010011 : VALUE=19'b0000000_100000100000;
      15'b011_111000010100 : VALUE=19'b0000000_100000011111;
      15'b011_111000010101 : VALUE=19'b0000000_100000011111;
      15'b011_111000010110 : VALUE=19'b0000000_100000011111;
      15'b011_111000010111 : VALUE=19'b0000000_100000011111;
      15'b011_111000011000 : VALUE=19'b0000000_100000011111;
      15'b011_111000011001 : VALUE=19'b0000000_100000011111;
      15'b011_111000011010 : VALUE=19'b0000000_100000011111;
      15'b011_111000011011 : VALUE=19'b0000000_100000011111;
      15'b011_111000011100 : VALUE=19'b0000000_100000011111;
      15'b011_111000011101 : VALUE=19'b0000000_100000011111;
      15'b011_111000011110 : VALUE=19'b0000000_100000011111;
      15'b011_111000011111 : VALUE=19'b0000000_100000011111;
      15'b011_111000100000 : VALUE=19'b0000000_100000011111;
      15'b011_111000100001 : VALUE=19'b0000000_100000011111;
      15'b011_111000100010 : VALUE=19'b0000000_100000011111;
      15'b011_111000100011 : VALUE=19'b0000000_100000011110;
      15'b011_111000100100 : VALUE=19'b0000000_100000011110;
      15'b011_111000100101 : VALUE=19'b0000000_100000011110;
      15'b011_111000100110 : VALUE=19'b0000000_100000011110;
      15'b011_111000100111 : VALUE=19'b0000000_100000011110;
      15'b011_111000101000 : VALUE=19'b0000000_100000011110;
      15'b011_111000101001 : VALUE=19'b0000000_100000011110;
      15'b011_111000101010 : VALUE=19'b0000000_100000011110;
      15'b011_111000101011 : VALUE=19'b0000000_100000011110;
      15'b011_111000101100 : VALUE=19'b0000000_100000011110;
      15'b011_111000101101 : VALUE=19'b0000000_100000011110;
      15'b011_111000101110 : VALUE=19'b0000000_100000011110;
      15'b011_111000101111 : VALUE=19'b0000000_100000011110;
      15'b011_111000110000 : VALUE=19'b0000000_100000011110;
      15'b011_111000110001 : VALUE=19'b0000000_100000011110;
      15'b011_111000110010 : VALUE=19'b0000000_100000011110;
      15'b011_111000110011 : VALUE=19'b0000000_100000011101;
      15'b011_111000110100 : VALUE=19'b0000000_100000011101;
      15'b011_111000110101 : VALUE=19'b0000000_100000011101;
      15'b011_111000110110 : VALUE=19'b0000000_100000011101;
      15'b011_111000110111 : VALUE=19'b0000000_100000011101;
      15'b011_111000111000 : VALUE=19'b0000000_100000011101;
      15'b011_111000111001 : VALUE=19'b0000000_100000011101;
      15'b011_111000111010 : VALUE=19'b0000000_100000011101;
      15'b011_111000111011 : VALUE=19'b0000000_100000011101;
      15'b011_111000111100 : VALUE=19'b0000000_100000011101;
      15'b011_111000111101 : VALUE=19'b0000000_100000011101;
      15'b011_111000111110 : VALUE=19'b0000000_100000011101;
      15'b011_111000111111 : VALUE=19'b0000000_100000011101;
      15'b011_111001000000 : VALUE=19'b0000000_100000011101;
      15'b011_111001000001 : VALUE=19'b0000000_100000011101;
      15'b011_111001000010 : VALUE=19'b0000000_100000011100;
      15'b011_111001000011 : VALUE=19'b0000000_100000011100;
      15'b011_111001000100 : VALUE=19'b0000000_100000011100;
      15'b011_111001000101 : VALUE=19'b0000000_100000011100;
      15'b011_111001000110 : VALUE=19'b0000000_100000011100;
      15'b011_111001000111 : VALUE=19'b0000000_100000011100;
      15'b011_111001001000 : VALUE=19'b0000000_100000011100;
      15'b011_111001001001 : VALUE=19'b0000000_100000011100;
      15'b011_111001001010 : VALUE=19'b0000000_100000011100;
      15'b011_111001001011 : VALUE=19'b0000000_100000011100;
      15'b011_111001001100 : VALUE=19'b0000000_100000011100;
      15'b011_111001001101 : VALUE=19'b0000000_100000011100;
      15'b011_111001001110 : VALUE=19'b0000000_100000011100;
      15'b011_111001001111 : VALUE=19'b0000000_100000011100;
      15'b011_111001010000 : VALUE=19'b0000000_100000011100;
      15'b011_111001010001 : VALUE=19'b0000000_100000011011;
      15'b011_111001010010 : VALUE=19'b0000000_100000011011;
      15'b011_111001010011 : VALUE=19'b0000000_100000011011;
      15'b011_111001010100 : VALUE=19'b0000000_100000011011;
      15'b011_111001010101 : VALUE=19'b0000000_100000011011;
      15'b011_111001010110 : VALUE=19'b0000000_100000011011;
      15'b011_111001010111 : VALUE=19'b0000000_100000011011;
      15'b011_111001011000 : VALUE=19'b0000000_100000011011;
      15'b011_111001011001 : VALUE=19'b0000000_100000011011;
      15'b011_111001011010 : VALUE=19'b0000000_100000011011;
      15'b011_111001011011 : VALUE=19'b0000000_100000011011;
      15'b011_111001011100 : VALUE=19'b0000000_100000011011;
      15'b011_111001011101 : VALUE=19'b0000000_100000011011;
      15'b011_111001011110 : VALUE=19'b0000000_100000011011;
      15'b011_111001011111 : VALUE=19'b0000000_100000011011;
      15'b011_111001100000 : VALUE=19'b0000000_100000011011;
      15'b011_111001100001 : VALUE=19'b0000000_100000011010;
      15'b011_111001100010 : VALUE=19'b0000000_100000011010;
      15'b011_111001100011 : VALUE=19'b0000000_100000011010;
      15'b011_111001100100 : VALUE=19'b0000000_100000011010;
      15'b011_111001100101 : VALUE=19'b0000000_100000011010;
      15'b011_111001100110 : VALUE=19'b0000000_100000011010;
      15'b011_111001100111 : VALUE=19'b0000000_100000011010;
      15'b011_111001101000 : VALUE=19'b0000000_100000011010;
      15'b011_111001101001 : VALUE=19'b0000000_100000011010;
      15'b011_111001101010 : VALUE=19'b0000000_100000011010;
      15'b011_111001101011 : VALUE=19'b0000000_100000011010;
      15'b011_111001101100 : VALUE=19'b0000000_100000011010;
      15'b011_111001101101 : VALUE=19'b0000000_100000011010;
      15'b011_111001101110 : VALUE=19'b0000000_100000011010;
      15'b011_111001101111 : VALUE=19'b0000000_100000011010;
      15'b011_111001110000 : VALUE=19'b0000000_100000011001;
      15'b011_111001110001 : VALUE=19'b0000000_100000011001;
      15'b011_111001110010 : VALUE=19'b0000000_100000011001;
      15'b011_111001110011 : VALUE=19'b0000000_100000011001;
      15'b011_111001110100 : VALUE=19'b0000000_100000011001;
      15'b011_111001110101 : VALUE=19'b0000000_100000011001;
      15'b011_111001110110 : VALUE=19'b0000000_100000011001;
      15'b011_111001110111 : VALUE=19'b0000000_100000011001;
      15'b011_111001111000 : VALUE=19'b0000000_100000011001;
      15'b011_111001111001 : VALUE=19'b0000000_100000011001;
      15'b011_111001111010 : VALUE=19'b0000000_100000011001;
      15'b011_111001111011 : VALUE=19'b0000000_100000011001;
      15'b011_111001111100 : VALUE=19'b0000000_100000011001;
      15'b011_111001111101 : VALUE=19'b0000000_100000011001;
      15'b011_111001111110 : VALUE=19'b0000000_100000011001;
      15'b011_111001111111 : VALUE=19'b0000000_100000011000;
      15'b011_111010000000 : VALUE=19'b0000000_100000011000;
      15'b011_111010000001 : VALUE=19'b0000000_100000011000;
      15'b011_111010000010 : VALUE=19'b0000000_100000011000;
      15'b011_111010000011 : VALUE=19'b0000000_100000011000;
      15'b011_111010000100 : VALUE=19'b0000000_100000011000;
      15'b011_111010000101 : VALUE=19'b0000000_100000011000;
      15'b011_111010000110 : VALUE=19'b0000000_100000011000;
      15'b011_111010000111 : VALUE=19'b0000000_100000011000;
      15'b011_111010001000 : VALUE=19'b0000000_100000011000;
      15'b011_111010001001 : VALUE=19'b0000000_100000011000;
      15'b011_111010001010 : VALUE=19'b0000000_100000011000;
      15'b011_111010001011 : VALUE=19'b0000000_100000011000;
      15'b011_111010001100 : VALUE=19'b0000000_100000011000;
      15'b011_111010001101 : VALUE=19'b0000000_100000011000;
      15'b011_111010001110 : VALUE=19'b0000000_100000011000;
      15'b011_111010001111 : VALUE=19'b0000000_100000010111;
      15'b011_111010010000 : VALUE=19'b0000000_100000010111;
      15'b011_111010010001 : VALUE=19'b0000000_100000010111;
      15'b011_111010010010 : VALUE=19'b0000000_100000010111;
      15'b011_111010010011 : VALUE=19'b0000000_100000010111;
      15'b011_111010010100 : VALUE=19'b0000000_100000010111;
      15'b011_111010010101 : VALUE=19'b0000000_100000010111;
      15'b011_111010010110 : VALUE=19'b0000000_100000010111;
      15'b011_111010010111 : VALUE=19'b0000000_100000010111;
      15'b011_111010011000 : VALUE=19'b0000000_100000010111;
      15'b011_111010011001 : VALUE=19'b0000000_100000010111;
      15'b011_111010011010 : VALUE=19'b0000000_100000010111;
      15'b011_111010011011 : VALUE=19'b0000000_100000010111;
      15'b011_111010011100 : VALUE=19'b0000000_100000010111;
      15'b011_111010011101 : VALUE=19'b0000000_100000010111;
      15'b011_111010011110 : VALUE=19'b0000000_100000010110;
      15'b011_111010011111 : VALUE=19'b0000000_100000010110;
      15'b011_111010100000 : VALUE=19'b0000000_100000010110;
      15'b011_111010100001 : VALUE=19'b0000000_100000010110;
      15'b011_111010100010 : VALUE=19'b0000000_100000010110;
      15'b011_111010100011 : VALUE=19'b0000000_100000010110;
      15'b011_111010100100 : VALUE=19'b0000000_100000010110;
      15'b011_111010100101 : VALUE=19'b0000000_100000010110;
      15'b011_111010100110 : VALUE=19'b0000000_100000010110;
      15'b011_111010100111 : VALUE=19'b0000000_100000010110;
      15'b011_111010101000 : VALUE=19'b0000000_100000010110;
      15'b011_111010101001 : VALUE=19'b0000000_100000010110;
      15'b011_111010101010 : VALUE=19'b0000000_100000010110;
      15'b011_111010101011 : VALUE=19'b0000000_100000010110;
      15'b011_111010101100 : VALUE=19'b0000000_100000010110;
      15'b011_111010101101 : VALUE=19'b0000000_100000010110;
      15'b011_111010101110 : VALUE=19'b0000000_100000010101;
      15'b011_111010101111 : VALUE=19'b0000000_100000010101;
      15'b011_111010110000 : VALUE=19'b0000000_100000010101;
      15'b011_111010110001 : VALUE=19'b0000000_100000010101;
      15'b011_111010110010 : VALUE=19'b0000000_100000010101;
      15'b011_111010110011 : VALUE=19'b0000000_100000010101;
      15'b011_111010110100 : VALUE=19'b0000000_100000010101;
      15'b011_111010110101 : VALUE=19'b0000000_100000010101;
      15'b011_111010110110 : VALUE=19'b0000000_100000010101;
      15'b011_111010110111 : VALUE=19'b0000000_100000010101;
      15'b011_111010111000 : VALUE=19'b0000000_100000010101;
      15'b011_111010111001 : VALUE=19'b0000000_100000010101;
      15'b011_111010111010 : VALUE=19'b0000000_100000010101;
      15'b011_111010111011 : VALUE=19'b0000000_100000010101;
      15'b011_111010111100 : VALUE=19'b0000000_100000010101;
      15'b011_111010111101 : VALUE=19'b0000000_100000010100;
      15'b011_111010111110 : VALUE=19'b0000000_100000010100;
      15'b011_111010111111 : VALUE=19'b0000000_100000010100;
      15'b011_111011000000 : VALUE=19'b0000000_100000010100;
      15'b011_111011000001 : VALUE=19'b0000000_100000010100;
      15'b011_111011000010 : VALUE=19'b0000000_100000010100;
      15'b011_111011000011 : VALUE=19'b0000000_100000010100;
      15'b011_111011000100 : VALUE=19'b0000000_100000010100;
      15'b011_111011000101 : VALUE=19'b0000000_100000010100;
      15'b011_111011000110 : VALUE=19'b0000000_100000010100;
      15'b011_111011000111 : VALUE=19'b0000000_100000010100;
      15'b011_111011001000 : VALUE=19'b0000000_100000010100;
      15'b011_111011001001 : VALUE=19'b0000000_100000010100;
      15'b011_111011001010 : VALUE=19'b0000000_100000010100;
      15'b011_111011001011 : VALUE=19'b0000000_100000010100;
      15'b011_111011001100 : VALUE=19'b0000000_100000010100;
      15'b011_111011001101 : VALUE=19'b0000000_100000010011;
      15'b011_111011001110 : VALUE=19'b0000000_100000010011;
      15'b011_111011001111 : VALUE=19'b0000000_100000010011;
      15'b011_111011010000 : VALUE=19'b0000000_100000010011;
      15'b011_111011010001 : VALUE=19'b0000000_100000010011;
      15'b011_111011010010 : VALUE=19'b0000000_100000010011;
      15'b011_111011010011 : VALUE=19'b0000000_100000010011;
      15'b011_111011010100 : VALUE=19'b0000000_100000010011;
      15'b011_111011010101 : VALUE=19'b0000000_100000010011;
      15'b011_111011010110 : VALUE=19'b0000000_100000010011;
      15'b011_111011010111 : VALUE=19'b0000000_100000010011;
      15'b011_111011011000 : VALUE=19'b0000000_100000010011;
      15'b011_111011011001 : VALUE=19'b0000000_100000010011;
      15'b011_111011011010 : VALUE=19'b0000000_100000010011;
      15'b011_111011011011 : VALUE=19'b0000000_100000010011;
      15'b011_111011011100 : VALUE=19'b0000000_100000010010;
      15'b011_111011011101 : VALUE=19'b0000000_100000010010;
      15'b011_111011011110 : VALUE=19'b0000000_100000010010;
      15'b011_111011011111 : VALUE=19'b0000000_100000010010;
      15'b011_111011100000 : VALUE=19'b0000000_100000010010;
      15'b011_111011100001 : VALUE=19'b0000000_100000010010;
      15'b011_111011100010 : VALUE=19'b0000000_100000010010;
      15'b011_111011100011 : VALUE=19'b0000000_100000010010;
      15'b011_111011100100 : VALUE=19'b0000000_100000010010;
      15'b011_111011100101 : VALUE=19'b0000000_100000010010;
      15'b011_111011100110 : VALUE=19'b0000000_100000010010;
      15'b011_111011100111 : VALUE=19'b0000000_100000010010;
      15'b011_111011101000 : VALUE=19'b0000000_100000010010;
      15'b011_111011101001 : VALUE=19'b0000000_100000010010;
      15'b011_111011101010 : VALUE=19'b0000000_100000010010;
      15'b011_111011101011 : VALUE=19'b0000000_100000010010;
      15'b011_111011101100 : VALUE=19'b0000000_100000010001;
      15'b011_111011101101 : VALUE=19'b0000000_100000010001;
      15'b011_111011101110 : VALUE=19'b0000000_100000010001;
      15'b011_111011101111 : VALUE=19'b0000000_100000010001;
      15'b011_111011110000 : VALUE=19'b0000000_100000010001;
      15'b011_111011110001 : VALUE=19'b0000000_100000010001;
      15'b011_111011110010 : VALUE=19'b0000000_100000010001;
      15'b011_111011110011 : VALUE=19'b0000000_100000010001;
      15'b011_111011110100 : VALUE=19'b0000000_100000010001;
      15'b011_111011110101 : VALUE=19'b0000000_100000010001;
      15'b011_111011110110 : VALUE=19'b0000000_100000010001;
      15'b011_111011110111 : VALUE=19'b0000000_100000010001;
      15'b011_111011111000 : VALUE=19'b0000000_100000010001;
      15'b011_111011111001 : VALUE=19'b0000000_100000010001;
      15'b011_111011111010 : VALUE=19'b0000000_100000010001;
      15'b011_111011111011 : VALUE=19'b0000000_100000010001;
      15'b011_111011111100 : VALUE=19'b0000000_100000010000;
      15'b011_111011111101 : VALUE=19'b0000000_100000010000;
      15'b011_111011111110 : VALUE=19'b0000000_100000010000;
      15'b011_111011111111 : VALUE=19'b0000000_100000010000;
      15'b011_111100000000 : VALUE=19'b0000000_100000010000;
      15'b011_111100000001 : VALUE=19'b0000000_100000010000;
      15'b011_111100000010 : VALUE=19'b0000000_100000010000;
      15'b011_111100000011 : VALUE=19'b0000000_100000010000;
      15'b011_111100000100 : VALUE=19'b0000000_100000010000;
      15'b011_111100000101 : VALUE=19'b0000000_100000010000;
      15'b011_111100000110 : VALUE=19'b0000000_100000010000;
      15'b011_111100000111 : VALUE=19'b0000000_100000010000;
      15'b011_111100001000 : VALUE=19'b0000000_100000010000;
      15'b011_111100001001 : VALUE=19'b0000000_100000010000;
      15'b011_111100001010 : VALUE=19'b0000000_100000010000;
      15'b011_111100001011 : VALUE=19'b0000000_100000001111;
      15'b011_111100001100 : VALUE=19'b0000000_100000001111;
      15'b011_111100001101 : VALUE=19'b0000000_100000001111;
      15'b011_111100001110 : VALUE=19'b0000000_100000001111;
      15'b011_111100001111 : VALUE=19'b0000000_100000001111;
      15'b011_111100010000 : VALUE=19'b0000000_100000001111;
      15'b011_111100010001 : VALUE=19'b0000000_100000001111;
      15'b011_111100010010 : VALUE=19'b0000000_100000001111;
      15'b011_111100010011 : VALUE=19'b0000000_100000001111;
      15'b011_111100010100 : VALUE=19'b0000000_100000001111;
      15'b011_111100010101 : VALUE=19'b0000000_100000001111;
      15'b011_111100010110 : VALUE=19'b0000000_100000001111;
      15'b011_111100010111 : VALUE=19'b0000000_100000001111;
      15'b011_111100011000 : VALUE=19'b0000000_100000001111;
      15'b011_111100011001 : VALUE=19'b0000000_100000001111;
      15'b011_111100011010 : VALUE=19'b0000000_100000001111;
      15'b011_111100011011 : VALUE=19'b0000000_100000001110;
      15'b011_111100011100 : VALUE=19'b0000000_100000001110;
      15'b011_111100011101 : VALUE=19'b0000000_100000001110;
      15'b011_111100011110 : VALUE=19'b0000000_100000001110;
      15'b011_111100011111 : VALUE=19'b0000000_100000001110;
      15'b011_111100100000 : VALUE=19'b0000000_100000001110;
      15'b011_111100100001 : VALUE=19'b0000000_100000001110;
      15'b011_111100100010 : VALUE=19'b0000000_100000001110;
      15'b011_111100100011 : VALUE=19'b0000000_100000001110;
      15'b011_111100100100 : VALUE=19'b0000000_100000001110;
      15'b011_111100100101 : VALUE=19'b0000000_100000001110;
      15'b011_111100100110 : VALUE=19'b0000000_100000001110;
      15'b011_111100100111 : VALUE=19'b0000000_100000001110;
      15'b011_111100101000 : VALUE=19'b0000000_100000001110;
      15'b011_111100101001 : VALUE=19'b0000000_100000001110;
      15'b011_111100101010 : VALUE=19'b0000000_100000001110;
      15'b011_111100101011 : VALUE=19'b0000000_100000001101;
      15'b011_111100101100 : VALUE=19'b0000000_100000001101;
      15'b011_111100101101 : VALUE=19'b0000000_100000001101;
      15'b011_111100101110 : VALUE=19'b0000000_100000001101;
      15'b011_111100101111 : VALUE=19'b0000000_100000001101;
      15'b011_111100110000 : VALUE=19'b0000000_100000001101;
      15'b011_111100110001 : VALUE=19'b0000000_100000001101;
      15'b011_111100110010 : VALUE=19'b0000000_100000001101;
      15'b011_111100110011 : VALUE=19'b0000000_100000001101;
      15'b011_111100110100 : VALUE=19'b0000000_100000001101;
      15'b011_111100110101 : VALUE=19'b0000000_100000001101;
      15'b011_111100110110 : VALUE=19'b0000000_100000001101;
      15'b011_111100110111 : VALUE=19'b0000000_100000001101;
      15'b011_111100111000 : VALUE=19'b0000000_100000001101;
      15'b011_111100111001 : VALUE=19'b0000000_100000001101;
      15'b011_111100111010 : VALUE=19'b0000000_100000001100;
      15'b011_111100111011 : VALUE=19'b0000000_100000001100;
      15'b011_111100111100 : VALUE=19'b0000000_100000001100;
      15'b011_111100111101 : VALUE=19'b0000000_100000001100;
      15'b011_111100111110 : VALUE=19'b0000000_100000001100;
      15'b011_111100111111 : VALUE=19'b0000000_100000001100;
      15'b011_111101000000 : VALUE=19'b0000000_100000001100;
      15'b011_111101000001 : VALUE=19'b0000000_100000001100;
      15'b011_111101000010 : VALUE=19'b0000000_100000001100;
      15'b011_111101000011 : VALUE=19'b0000000_100000001100;
      15'b011_111101000100 : VALUE=19'b0000000_100000001100;
      15'b011_111101000101 : VALUE=19'b0000000_100000001100;
      15'b011_111101000110 : VALUE=19'b0000000_100000001100;
      15'b011_111101000111 : VALUE=19'b0000000_100000001100;
      15'b011_111101001000 : VALUE=19'b0000000_100000001100;
      15'b011_111101001001 : VALUE=19'b0000000_100000001100;
      15'b011_111101001010 : VALUE=19'b0000000_100000001011;
      15'b011_111101001011 : VALUE=19'b0000000_100000001011;
      15'b011_111101001100 : VALUE=19'b0000000_100000001011;
      15'b011_111101001101 : VALUE=19'b0000000_100000001011;
      15'b011_111101001110 : VALUE=19'b0000000_100000001011;
      15'b011_111101001111 : VALUE=19'b0000000_100000001011;
      15'b011_111101010000 : VALUE=19'b0000000_100000001011;
      15'b011_111101010001 : VALUE=19'b0000000_100000001011;
      15'b011_111101010010 : VALUE=19'b0000000_100000001011;
      15'b011_111101010011 : VALUE=19'b0000000_100000001011;
      15'b011_111101010100 : VALUE=19'b0000000_100000001011;
      15'b011_111101010101 : VALUE=19'b0000000_100000001011;
      15'b011_111101010110 : VALUE=19'b0000000_100000001011;
      15'b011_111101010111 : VALUE=19'b0000000_100000001011;
      15'b011_111101011000 : VALUE=19'b0000000_100000001011;
      15'b011_111101011001 : VALUE=19'b0000000_100000001011;
      15'b011_111101011010 : VALUE=19'b0000000_100000001010;
      15'b011_111101011011 : VALUE=19'b0000000_100000001010;
      15'b011_111101011100 : VALUE=19'b0000000_100000001010;
      15'b011_111101011101 : VALUE=19'b0000000_100000001010;
      15'b011_111101011110 : VALUE=19'b0000000_100000001010;
      15'b011_111101011111 : VALUE=19'b0000000_100000001010;
      15'b011_111101100000 : VALUE=19'b0000000_100000001010;
      15'b011_111101100001 : VALUE=19'b0000000_100000001010;
      15'b011_111101100010 : VALUE=19'b0000000_100000001010;
      15'b011_111101100011 : VALUE=19'b0000000_100000001010;
      15'b011_111101100100 : VALUE=19'b0000000_100000001010;
      15'b011_111101100101 : VALUE=19'b0000000_100000001010;
      15'b011_111101100110 : VALUE=19'b0000000_100000001010;
      15'b011_111101100111 : VALUE=19'b0000000_100000001010;
      15'b011_111101101000 : VALUE=19'b0000000_100000001010;
      15'b011_111101101001 : VALUE=19'b0000000_100000001010;
      15'b011_111101101010 : VALUE=19'b0000000_100000001001;
      15'b011_111101101011 : VALUE=19'b0000000_100000001001;
      15'b011_111101101100 : VALUE=19'b0000000_100000001001;
      15'b011_111101101101 : VALUE=19'b0000000_100000001001;
      15'b011_111101101110 : VALUE=19'b0000000_100000001001;
      15'b011_111101101111 : VALUE=19'b0000000_100000001001;
      15'b011_111101110000 : VALUE=19'b0000000_100000001001;
      15'b011_111101110001 : VALUE=19'b0000000_100000001001;
      15'b011_111101110010 : VALUE=19'b0000000_100000001001;
      15'b011_111101110011 : VALUE=19'b0000000_100000001001;
      15'b011_111101110100 : VALUE=19'b0000000_100000001001;
      15'b011_111101110101 : VALUE=19'b0000000_100000001001;
      15'b011_111101110110 : VALUE=19'b0000000_100000001001;
      15'b011_111101110111 : VALUE=19'b0000000_100000001001;
      15'b011_111101111000 : VALUE=19'b0000000_100000001001;
      15'b011_111101111001 : VALUE=19'b0000000_100000001000;
      15'b011_111101111010 : VALUE=19'b0000000_100000001000;
      15'b011_111101111011 : VALUE=19'b0000000_100000001000;
      15'b011_111101111100 : VALUE=19'b0000000_100000001000;
      15'b011_111101111101 : VALUE=19'b0000000_100000001000;
      15'b011_111101111110 : VALUE=19'b0000000_100000001000;
      15'b011_111101111111 : VALUE=19'b0000000_100000001000;
      15'b011_111110000000 : VALUE=19'b0000000_100000001000;
      15'b011_111110000001 : VALUE=19'b0000000_100000001000;
      15'b011_111110000010 : VALUE=19'b0000000_100000001000;
      15'b011_111110000011 : VALUE=19'b0000000_100000001000;
      15'b011_111110000100 : VALUE=19'b0000000_100000001000;
      15'b011_111110000101 : VALUE=19'b0000000_100000001000;
      15'b011_111110000110 : VALUE=19'b0000000_100000001000;
      15'b011_111110000111 : VALUE=19'b0000000_100000001000;
      15'b011_111110001000 : VALUE=19'b0000000_100000001000;
      15'b011_111110001001 : VALUE=19'b0000000_100000000111;
      15'b011_111110001010 : VALUE=19'b0000000_100000000111;
      15'b011_111110001011 : VALUE=19'b0000000_100000000111;
      15'b011_111110001100 : VALUE=19'b0000000_100000000111;
      15'b011_111110001101 : VALUE=19'b0000000_100000000111;
      15'b011_111110001110 : VALUE=19'b0000000_100000000111;
      15'b011_111110001111 : VALUE=19'b0000000_100000000111;
      15'b011_111110010000 : VALUE=19'b0000000_100000000111;
      15'b011_111110010001 : VALUE=19'b0000000_100000000111;
      15'b011_111110010010 : VALUE=19'b0000000_100000000111;
      15'b011_111110010011 : VALUE=19'b0000000_100000000111;
      15'b011_111110010100 : VALUE=19'b0000000_100000000111;
      15'b011_111110010101 : VALUE=19'b0000000_100000000111;
      15'b011_111110010110 : VALUE=19'b0000000_100000000111;
      15'b011_111110010111 : VALUE=19'b0000000_100000000111;
      15'b011_111110011000 : VALUE=19'b0000000_100000000111;
      15'b011_111110011001 : VALUE=19'b0000000_100000000110;
      15'b011_111110011010 : VALUE=19'b0000000_100000000110;
      15'b011_111110011011 : VALUE=19'b0000000_100000000110;
      15'b011_111110011100 : VALUE=19'b0000000_100000000110;
      15'b011_111110011101 : VALUE=19'b0000000_100000000110;
      15'b011_111110011110 : VALUE=19'b0000000_100000000110;
      15'b011_111110011111 : VALUE=19'b0000000_100000000110;
      15'b011_111110100000 : VALUE=19'b0000000_100000000110;
      15'b011_111110100001 : VALUE=19'b0000000_100000000110;
      15'b011_111110100010 : VALUE=19'b0000000_100000000110;
      15'b011_111110100011 : VALUE=19'b0000000_100000000110;
      15'b011_111110100100 : VALUE=19'b0000000_100000000110;
      15'b011_111110100101 : VALUE=19'b0000000_100000000110;
      15'b011_111110100110 : VALUE=19'b0000000_100000000110;
      15'b011_111110100111 : VALUE=19'b0000000_100000000110;
      15'b011_111110101000 : VALUE=19'b0000000_100000000110;
      15'b011_111110101001 : VALUE=19'b0000000_100000000101;
      15'b011_111110101010 : VALUE=19'b0000000_100000000101;
      15'b011_111110101011 : VALUE=19'b0000000_100000000101;
      15'b011_111110101100 : VALUE=19'b0000000_100000000101;
      15'b011_111110101101 : VALUE=19'b0000000_100000000101;
      15'b011_111110101110 : VALUE=19'b0000000_100000000101;
      15'b011_111110101111 : VALUE=19'b0000000_100000000101;
      15'b011_111110110000 : VALUE=19'b0000000_100000000101;
      15'b011_111110110001 : VALUE=19'b0000000_100000000101;
      15'b011_111110110010 : VALUE=19'b0000000_100000000101;
      15'b011_111110110011 : VALUE=19'b0000000_100000000101;
      15'b011_111110110100 : VALUE=19'b0000000_100000000101;
      15'b011_111110110101 : VALUE=19'b0000000_100000000101;
      15'b011_111110110110 : VALUE=19'b0000000_100000000101;
      15'b011_111110110111 : VALUE=19'b0000000_100000000101;
      15'b011_111110111000 : VALUE=19'b0000000_100000000101;
      15'b011_111110111001 : VALUE=19'b0000000_100000000100;
      15'b011_111110111010 : VALUE=19'b0000000_100000000100;
      15'b011_111110111011 : VALUE=19'b0000000_100000000100;
      15'b011_111110111100 : VALUE=19'b0000000_100000000100;
      15'b011_111110111101 : VALUE=19'b0000000_100000000100;
      15'b011_111110111110 : VALUE=19'b0000000_100000000100;
      15'b011_111110111111 : VALUE=19'b0000000_100000000100;
      15'b011_111111000000 : VALUE=19'b0000000_100000000100;
      15'b011_111111000001 : VALUE=19'b0000000_100000000100;
      15'b011_111111000010 : VALUE=19'b0000000_100000000100;
      15'b011_111111000011 : VALUE=19'b0000000_100000000100;
      15'b011_111111000100 : VALUE=19'b0000000_100000000100;
      15'b011_111111000101 : VALUE=19'b0000000_100000000100;
      15'b011_111111000110 : VALUE=19'b0000000_100000000100;
      15'b011_111111000111 : VALUE=19'b0000000_100000000100;
      15'b011_111111001000 : VALUE=19'b0000000_100000000100;
      15'b011_111111001001 : VALUE=19'b0000000_100000000011;
      15'b011_111111001010 : VALUE=19'b0000000_100000000011;
      15'b011_111111001011 : VALUE=19'b0000000_100000000011;
      15'b011_111111001100 : VALUE=19'b0000000_100000000011;
      15'b011_111111001101 : VALUE=19'b0000000_100000000011;
      15'b011_111111001110 : VALUE=19'b0000000_100000000011;
      15'b011_111111001111 : VALUE=19'b0000000_100000000011;
      15'b011_111111010000 : VALUE=19'b0000000_100000000011;
      15'b011_111111010001 : VALUE=19'b0000000_100000000011;
      15'b011_111111010010 : VALUE=19'b0000000_100000000011;
      15'b011_111111010011 : VALUE=19'b0000000_100000000011;
      15'b011_111111010100 : VALUE=19'b0000000_100000000011;
      15'b011_111111010101 : VALUE=19'b0000000_100000000011;
      15'b011_111111010110 : VALUE=19'b0000000_100000000011;
      15'b011_111111010111 : VALUE=19'b0000000_100000000011;
      15'b011_111111011000 : VALUE=19'b0000000_100000000011;
      15'b011_111111011001 : VALUE=19'b0000000_100000000010;
      15'b011_111111011010 : VALUE=19'b0000000_100000000010;
      15'b011_111111011011 : VALUE=19'b0000000_100000000010;
      15'b011_111111011100 : VALUE=19'b0000000_100000000010;
      15'b011_111111011101 : VALUE=19'b0000000_100000000010;
      15'b011_111111011110 : VALUE=19'b0000000_100000000010;
      15'b011_111111011111 : VALUE=19'b0000000_100000000010;
      15'b011_111111100000 : VALUE=19'b0000000_100000000010;
      15'b011_111111100001 : VALUE=19'b0000000_100000000010;
      15'b011_111111100010 : VALUE=19'b0000000_100000000010;
      15'b011_111111100011 : VALUE=19'b0000000_100000000010;
      15'b011_111111100100 : VALUE=19'b0000000_100000000010;
      15'b011_111111100101 : VALUE=19'b0000000_100000000010;
      15'b011_111111100110 : VALUE=19'b0000000_100000000010;
      15'b011_111111100111 : VALUE=19'b0000000_100000000010;
      15'b011_111111101000 : VALUE=19'b0000000_100000000010;
      15'b011_111111101001 : VALUE=19'b0000000_100000000001;
      15'b011_111111101010 : VALUE=19'b0000000_100000000001;
      15'b011_111111101011 : VALUE=19'b0000000_100000000001;
      15'b011_111111101100 : VALUE=19'b0000000_100000000001;
      15'b011_111111101101 : VALUE=19'b0000000_100000000001;
      15'b011_111111101110 : VALUE=19'b0000000_100000000001;
      15'b011_111111101111 : VALUE=19'b0000000_100000000001;
      15'b011_111111110000 : VALUE=19'b0000000_100000000001;
      15'b011_111111110001 : VALUE=19'b0000000_100000000001;
      15'b011_111111110010 : VALUE=19'b0000000_100000000001;
      15'b011_111111110011 : VALUE=19'b0000000_100000000001;
      15'b011_111111110100 : VALUE=19'b0000000_100000000001;
      15'b011_111111110101 : VALUE=19'b0000000_100000000001;
      15'b011_111111110110 : VALUE=19'b0000000_100000000001;
      15'b011_111111110111 : VALUE=19'b0000000_100000000001;
      15'b011_111111111000 : VALUE=19'b0000000_100000000001;
      15'b011_111111111001 : VALUE=19'b0000000_100000000000;
      15'b011_111111111010 : VALUE=19'b0000000_100000000000;
      15'b011_111111111011 : VALUE=19'b0000000_100000000000;
      15'b011_111111111100 : VALUE=19'b0000000_100000000000;
      15'b011_111111111101 : VALUE=19'b0000000_100000000000;
      15'b011_111111111110 : VALUE=19'b0000000_100000000000;
      15'b011_111111111111 : VALUE=19'b0000000_100000000000;
    endcase
  end
endmodule
